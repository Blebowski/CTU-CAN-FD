--------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core
-- Copyright (C) 2015-2018
-- 
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
-- 
-- Project advisors: 
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
-- 
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Memory map for: CAN_Frame_format
-- This file is autogenerated, DO NOT EDIT!
--------------------------------------------------------------------------------

Library ieee;
use ieee.std_logic_1164.all;

package can_fd_frame_format is

  ------------------------------------------------------------------------------
  -- Common types
  ------------------------------------------------------------------------------
  type t_reg_type is (
    reg_none,
    reg_write_only,
    reg_read_only,
    reg_read_write,
    reg_read_write_once
  );

  type t_memory_reg is record
       address       : std_logic_vector(11 downto 0);
       size                                : integer;
       reg_type                         : t_reg_type;
       reset_val     : std_logic_vector(31 downto 0);
       is_implem     : std_logic_vector(31 downto 0);
  end record;


  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: CAN_FD_Frame_format
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant CAN_FD_FRAME_FORMAT_BLOCK    : std_logic_vector(3 downto 0) := x"0";

  constant FRAME_FORM_W_ADR          : std_logic_vector(11 downto 0) := x"000";
  constant IDENTIFIER_W_ADR          : std_logic_vector(11 downto 0) := x"004";
  constant TIMESTAMP_L_W_ADR         : std_logic_vector(11 downto 0) := x"008";
  constant TIMESTAMP_U_W_ADR         : std_logic_vector(11 downto 0) := x"00C";
  constant DATA_1_4_W_ADR            : std_logic_vector(11 downto 0) := x"010";
  constant DATA_5_8_W_ADR            : std_logic_vector(11 downto 0) := x"014";
  constant DATA_61_64_W_ADR          : std_logic_vector(11 downto 0) := x"04C";

  ------------------------------------------------------------------------------
  -- Register list
  ------------------------------------------------------------------------------

  type t_CAN_FD_Frame_format_list is array (0 to 6) of t_memory_reg;

  constant CAN_FD_Frame_format_list : t_CAN_FD_Frame_format_list :=(

    (address   => FRAME_FORM_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "00000000000000001111111011101111"),
    (address   => IDENTIFIER_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "00011111111111111111111111111111"),
    (address   => TIMESTAMP_L_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "11111111111111111111111111111111"),
    (address   => TIMESTAMP_U_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "11111111111111111111111111111111"),
    (address   => DATA_1_4_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "11111111111111111111111111111111"),
    (address   => DATA_5_8_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "11111111111111111111111111111111"),
    (address   => DATA_61_64_W_ADR,
     size      => 32,
     reg_type  => reg_none,
     reset_val => "00000000000000000000000000000000",
     is_implem => "11111111111111111111111111111111")
  );

  ------------------------------------------------------------------------------
  -- FRAME_FORM_W register
  --
  -- Frame format word with CAN frame metadata.
  ------------------------------------------------------------------------------
  constant DLC_L                  : natural := 0;
  constant DLC_H                  : natural := 3;
  constant RTR_IND                : natural := 5;
  constant IDE_IND                : natural := 6;
  constant FDF_IND                : natural := 7;
  constant BRS_IND                : natural := 9;
  constant ESI_RSV_IND           : natural := 10;
  constant RWCNT_L               : natural := 11;
  constant RWCNT_H               : natural := 15;

  -- "RTR" field enumerated values
  constant NO_RTR_FRAME       : std_logic := '0';
  constant RTR_FRAME          : std_logic := '1';

  -- "IDE" field enumerated values
  constant BASE               : std_logic := '0';
  constant EXTENDED           : std_logic := '1';

  -- "FDF" field enumerated values
  constant NORMAL_CAN         : std_logic := '0';
  constant FD_CAN             : std_logic := '1';

  -- "BRS" field enumerated values
  constant BR_NO_SHIFT        : std_logic := '0';
  constant BR_SHIFT           : std_logic := '1';

  -- "ESI_RSV" field enumerated values
  constant ESI_ERR_ACTIVE     : std_logic := '0';
  constant ESI_ERR_PASIVE     : std_logic := '1';

  -- FRAME_FORM_W register reset values

  ------------------------------------------------------------------------------
  -- IDENTIFIER_W register
  --
  -- CAN Identifier.
  ------------------------------------------------------------------------------
  constant IDENTIFIER_EXT_L       : natural := 0;
  constant IDENTIFIER_EXT_H      : natural := 17;
  constant IDENTIFIER_BASE_L     : natural := 18;
  constant IDENTIFIER_BASE_H     : natural := 28;

  -- IDENTIFIER_W register reset values

  ------------------------------------------------------------------------------
  -- TIMESTAMP_L_W register
  --
  ------------------------------------------------------------------------------
  constant TIME_STAMP_31_0_L      : natural := 0;
  constant TIME_STAMP_31_0_H     : natural := 31;

  -- TIMESTAMP_L_W register reset values

  ------------------------------------------------------------------------------
  -- TIMESTAMP_U_W register
  --
  ------------------------------------------------------------------------------
  constant TIMESTAMP_L_W_L        : natural := 0;
  constant TIMESTAMP_L_W_H       : natural := 31;

  -- TIMESTAMP_U_W register reset values

  ------------------------------------------------------------------------------
  -- DATA_1_4_W register
  --
  ------------------------------------------------------------------------------
  constant DATA_1_L               : natural := 0;
  constant DATA_1_H               : natural := 7;
  constant DATA_2_L               : natural := 8;
  constant DATA_2_H              : natural := 15;
  constant DATA_3_L              : natural := 16;
  constant DATA_3_H              : natural := 23;
  constant DATA_4_L              : natural := 24;
  constant DATA_4_H              : natural := 31;

  -- DATA_1_4_W register reset values

  ------------------------------------------------------------------------------
  -- DATA_5_8_W register
  --
  ------------------------------------------------------------------------------
  constant DATA_5_L               : natural := 0;
  constant DATA_5_H               : natural := 7;
  constant DATA_6_L               : natural := 8;
  constant DATA_6_H              : natural := 15;
  constant DATA_7_L              : natural := 16;
  constant DATA_7_H              : natural := 23;
  constant DATA_8_L              : natural := 24;
  constant DATA_8_H              : natural := 31;

  -- DATA_5_8_W register reset values

  ------------------------------------------------------------------------------
  -- DATA_61_64_W register
  --
  ------------------------------------------------------------------------------
  constant DATA_61_L              : natural := 0;
  constant DATA_61_H              : natural := 7;
  constant DATA_62_L              : natural := 8;
  constant DATA_62_H             : natural := 15;
  constant DATA_63_L             : natural := 16;
  constant DATA_63_H             : natural := 23;
  constant DATA_64_L             : natural := 24;
  constant DATA_64_H             : natural := 31;

  -- DATA_61_64_W register reset values

end package;
