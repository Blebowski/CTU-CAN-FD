--------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core
-- Copyright (C) 2015-2018
-- 
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
-- 
-- Project advisors: 
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
-- 
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- Memory map for: CAN_Registers
-- This file is autogenerated, DO NOT EDIT!
--------------------------------------------------------------------------------

Library ieee;
use ieee.std_logic_1164.all;

package can_fd_register_map is

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: Control_registers
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant CONTROL_REGISTERS_BLOCK      : std_logic_vector(3 downto 0) := x"0";

  constant DEVICE_ID_ADR             : std_logic_vector(11 downto 0) := x"000";
  constant VERSION_ADR               : std_logic_vector(11 downto 0) := x"002";
  constant MODE_ADR                  : std_logic_vector(11 downto 0) := x"004";
  constant COMMAND_ADR               : std_logic_vector(11 downto 0) := x"005";
  constant STATUS_ADR                : std_logic_vector(11 downto 0) := x"006";
  constant SETTINGS_ADR              : std_logic_vector(11 downto 0) := x"007";
  constant INT_STAT_ADR              : std_logic_vector(11 downto 0) := x"008";
  constant INT_ENA_SET_ADR           : std_logic_vector(11 downto 0) := x"00C";
  constant INT_ENA_CLR_ADR           : std_logic_vector(11 downto 0) := x"010";
  constant INT_MASK_SET_ADR          : std_logic_vector(11 downto 0) := x"014";
  constant INT_MASK_CLR_ADR          : std_logic_vector(11 downto 0) := x"018";
  constant BTR_ADR                   : std_logic_vector(11 downto 0) := x"01C";
  constant BTR_FD_ADR                : std_logic_vector(11 downto 0) := x"020";
  constant EWL_ADR                   : std_logic_vector(11 downto 0) := x"024";
  constant ERP_ADR                   : std_logic_vector(11 downto 0) := x"025";
  constant FAULT_STATE_ADR           : std_logic_vector(11 downto 0) := x"026";
  constant RXC_ADR                   : std_logic_vector(11 downto 0) := x"028";
  constant TXC_ADR                   : std_logic_vector(11 downto 0) := x"02A";
  constant ERR_NORM_ADR              : std_logic_vector(11 downto 0) := x"02C";
  constant ERR_FD_ADR                : std_logic_vector(11 downto 0) := x"02E";
  constant CTR_PRES_ADR              : std_logic_vector(11 downto 0) := x"030";
  constant FILTER_A_MASK_ADR         : std_logic_vector(11 downto 0) := x"034";
  constant FILTER_A_VAL_ADR          : std_logic_vector(11 downto 0) := x"038";
  constant FILTER_B_MASK_ADR         : std_logic_vector(11 downto 0) := x"03C";
  constant FILTER_B_VAL_ADR          : std_logic_vector(11 downto 0) := x"040";
  constant FILTER_C_MASK_ADR         : std_logic_vector(11 downto 0) := x"044";
  constant FILTER_C_VAL_ADR          : std_logic_vector(11 downto 0) := x"048";
  constant FILTER_RAN_LOW_ADR        : std_logic_vector(11 downto 0) := x"04C";
  constant FILTER_RAN_HIGH_ADR       : std_logic_vector(11 downto 0) := x"050";
  constant FILTER_CONTROL_ADR        : std_logic_vector(11 downto 0) := x"054";
  constant FILTER_STATUS_ADR         : std_logic_vector(11 downto 0) := x"056";
  constant RX_MEM_INFO_ADR           : std_logic_vector(11 downto 0) := x"058";
  constant RX_POINTERS_ADR           : std_logic_vector(11 downto 0) := x"05C";
  constant RX_STATUS_ADR             : std_logic_vector(11 downto 0) := x"060";
  constant RX_SETTINGS_ADR           : std_logic_vector(11 downto 0) := x"062";
  constant RX_DATA_ADR               : std_logic_vector(11 downto 0) := x"064";
  constant TX_STATUS_ADR             : std_logic_vector(11 downto 0) := x"068";
  constant TX_COMMAND_ADR            : std_logic_vector(11 downto 0) := x"06C";
  constant TX_PRIORITY_ADR           : std_logic_vector(11 downto 0) := x"070";
  constant ERR_CAPT_ADR              : std_logic_vector(11 downto 0) := x"074";
  constant ALC_ADR                   : std_logic_vector(11 downto 0) := x"075";
  constant TRV_DELAY_ADR             : std_logic_vector(11 downto 0) := x"078";
  constant SSP_CFG_ADR               : std_logic_vector(11 downto 0) := x"07A";
  constant RX_COUNTER_ADR            : std_logic_vector(11 downto 0) := x"07C";
  constant TX_COUNTER_ADR            : std_logic_vector(11 downto 0) := x"080";
  constant DEBUG_REGISTER_ADR        : std_logic_vector(11 downto 0) := x"084";
  constant YOLO_REG_ADR              : std_logic_vector(11 downto 0) := x"088";
  constant TIMESTAMP_LOW_ADR         : std_logic_vector(11 downto 0) := x"08C";
  constant TIMESTAMP_HIGH_ADR        : std_logic_vector(11 downto 0) := x"090";

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: TX_Buffer_1
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant TX_BUFFER_1_BLOCK            : std_logic_vector(3 downto 0) := x"1";

  constant TXTB1_DATA_1_ADR          : std_logic_vector(11 downto 0) := x"100";
  constant TXTB1_DATA_2_ADR          : std_logic_vector(11 downto 0) := x"104";
  constant TXTB1_DATA_20_ADR         : std_logic_vector(11 downto 0) := x"14C";

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: TX_Buffer_2
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant TX_BUFFER_2_BLOCK            : std_logic_vector(3 downto 0) := x"2";

  constant TXTB2_DATA_1_ADR          : std_logic_vector(11 downto 0) := x"200";
  constant TXTB2_DATA_2_ADR          : std_logic_vector(11 downto 0) := x"204";
  constant TXTB2_DATA_20_ADR         : std_logic_vector(11 downto 0) := x"24C";

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: TX_Buffer_3
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant TX_BUFFER_3_BLOCK            : std_logic_vector(3 downto 0) := x"3";

  constant TXTB3_DATA_1_ADR          : std_logic_vector(11 downto 0) := x"300";
  constant TXTB3_DATA_2_ADR          : std_logic_vector(11 downto 0) := x"304";
  constant TXTB3_DATA_20_ADR         : std_logic_vector(11 downto 0) := x"34C";

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: TX_Buffer_4
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant TX_BUFFER_4_BLOCK            : std_logic_vector(3 downto 0) := x"4";

  constant TXTB4_DATA_1_ADR          : std_logic_vector(11 downto 0) := x"400";
  constant TXTB4_DATA_2_ADR          : std_logic_vector(11 downto 0) := x"404";
  constant TXTB4_DATA_20_ADR         : std_logic_vector(11 downto 0) := x"44C";

  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  -- Address block: Event_Logger
  ------------------------------------------------------------------------------
  ------------------------------------------------------------------------------
  constant EVENT_LOGGER_BLOCK           : std_logic_vector(3 downto 0) := x"5";

  constant LOG_TRIG_CONFIG_ADR       : std_logic_vector(11 downto 0) := x"500";
  constant LOG_CAPT_CONFIG_ADR       : std_logic_vector(11 downto 0) := x"504";
  constant LOG_STATUS_ADR            : std_logic_vector(11 downto 0) := x"508";
  constant LOG_POINTERS_ADR          : std_logic_vector(11 downto 0) := x"50A";
  constant LOG_COMMAND_ADR           : std_logic_vector(11 downto 0) := x"50C";
  constant LOG_CAPT_EVENT_1_ADR      : std_logic_vector(11 downto 0) := x"510";
  constant LOG_CAPT_EVENT_2_ADR      : std_logic_vector(11 downto 0) := x"514";

  ------------------------------------------------------------------------------
  -- DEVICE_ID register
  --
  -- Register contains the identifer of CTU CAN FD IP Core. It can be used to de
  -- termine if CTU CAN FD IP Core is mapped correctly on its base address.
  ------------------------------------------------------------------------------
  constant DEVICE_ID_L            : natural := 0;
  constant DEVICE_ID_H           : natural := 15;

  -- "DEVICE_ID" field enumerated values
  constant CTU_CAN_FD_ID : std_logic_vector(15 downto 0) := x"CAFD";

  -- DEVICE_ID register reset values
  constant DEVICE_ID_RSTVAL : std_logic_vector(15 downto 0) := x"CAFD";

  ------------------------------------------------------------------------------
  -- VERSION register
  --
  -- Version register with IP Core version.
  ------------------------------------------------------------------------------
  constant VER_MINOR_L           : natural := 16;
  constant VER_MINOR_H           : natural := 23;
  constant VER_MAJOR_L           : natural := 24;
  constant VER_MAJOR_H           : natural := 31;

  -- VERSION register reset values

  ------------------------------------------------------------------------------
  -- MODE register
  --
  -- MODE register controls operating modes.
  ------------------------------------------------------------------------------
  constant RST_IND                : natural := 0;
  constant LOM_IND                : natural := 1;
  constant STM_IND                : natural := 2;
  constant AFM_IND                : natural := 3;
  constant FDE_IND                : natural := 4;
  constant RTRP_IND               : natural := 5;
  constant TSM_IND                : natural := 6;
  constant ACF_IND                : natural := 7;

  -- "FDE" field enumerated values
  constant FDE_DISABLE        : std_logic := '0';
  constant FDE_ENABLE         : std_logic := '1';

  -- "TSM" field enumerated values
  constant TSM_DISABLE        : std_logic := '0';
  constant TSM_ENABLE         : std_logic := '1';

  -- "RTRP" field enumerated values
  constant RTR_EXTRA          : std_logic := '0';
  constant RTR_STANDARD       : std_logic := '1';

  -- "ACF" field enumerated values
  constant ACF_DISABLED       : std_logic := '0';
  constant ACF_ENABLED        : std_logic := '1';

  -- "LOM" field enumerated values
  constant LOM_DISABLED       : std_logic := '0';
  constant LOM_ENABLED        : std_logic := '1';

  -- "STM" field enumerated values
  constant STM_DISABLED       : std_logic := '0';
  constant STM_ENABLED        : std_logic := '1';

  -- "AFM" field enumerated values
  constant AFM_DISABLED       : std_logic := '0';
  constant AFM_ENABLED        : std_logic := '1';

  -- MODE register reset values
  constant RST_RSTVAL         : std_logic := '0';
  constant FDE_RSTVAL         : std_logic := '1';
  constant TSM_RSTVAL         : std_logic := '0';
  constant RTRP_RSTVAL        : std_logic := '1';
  constant ACF_RSTVAL         : std_logic := '0';
  constant LOM_RSTVAL         : std_logic := '0';
  constant STM_RSTVAL         : std_logic := '0';
  constant AFM_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- COMMAND register
  --
  -- Writing logic 1 into each bit gives different command to the IP Core. After
  --  writing logic 1, logic 0 does not have to be written.
  ------------------------------------------------------------------------------
  constant ABT_IND                : natural := 9;
  constant RRB_IND               : natural := 10;
  constant CDO_IND               : natural := 11;
  constant ERCRST_IND            : natural := 12;
  constant RXFCRST_IND           : natural := 13;
  constant TXFCRST_IND           : natural := 14;

  -- COMMAND register reset values
  constant ABT_RSTVAL         : std_logic := '0';
  constant RRB_RSTVAL         : std_logic := '0';
  constant CDO_RSTVAL         : std_logic := '0';
  constant ERCRST_RSTVAL      : std_logic := '0';
  constant RXFCRST_RSTVAL     : std_logic := '0';
  constant TXFCRST_RSTVAL     : std_logic := '0';

  ------------------------------------------------------------------------------
  -- STATUS register
  --
  -- Register signals various states of CTU CAN FD IP Core. Logic 1 signals acti
  -- ve status/flag.
  ------------------------------------------------------------------------------
  constant RXNE_IND              : natural := 16;
  constant DOR_IND               : natural := 17;
  constant TXNF_IND              : natural := 18;
  constant EFT_IND               : natural := 19;
  constant RXS_IND               : natural := 20;
  constant TXS_IND               : natural := 21;
  constant EWL_IND               : natural := 22;
  constant IDLE_IND              : natural := 23;

  -- STATUS register reset values
  constant RXNE_RSTVAL        : std_logic := '0';
  constant TXNF_RSTVAL        : std_logic := '0';
  constant DOR_RSTVAL         : std_logic := '0';
  constant EFT_RSTVAL         : std_logic := '0';
  constant RXS_RSTVAL         : std_logic := '0';
  constant TXS_RSTVAL         : std_logic := '0';
  constant EWL_RSTVAL         : std_logic := '0';
  constant IDLE_RSTVAL        : std_logic := '1';

  ------------------------------------------------------------------------------
  -- SETTINGS register
  --
  -- This register enables the whole CAN FD Core, configures FD Type, Internal l
  -- oopback and retransmission options.
  ------------------------------------------------------------------------------
  constant RTRLE_IND             : natural := 24;
  constant RTRTH_L               : natural := 25;
  constant RTRTH_H               : natural := 28;
  constant ILBP_IND              : natural := 29;
  constant ENA_IND               : natural := 30;
  constant NISOFD_IND            : natural := 31;

  -- "RTRLE" field enumerated values
  constant RTRLE_DISABLED     : std_logic := '0';
  constant RTRLE_ENABLED      : std_logic := '1';

  -- "ILBP" field enumerated values
  constant INT_LOOP_DISABLED  : std_logic := '0';
  constant INT_LOOP_ENABLED   : std_logic := '1';

  -- "ENA" field enumerated values
  constant DISABLED           : std_logic := '0';
  constant ENABLED            : std_logic := '1';

  -- "NISOFD" field enumerated values
  constant ISO_FD             : std_logic := '0';
  constant NON_ISO_FD         : std_logic := '1';

  -- SETTINGS register reset values
  constant RTRLE_RSTVAL       : std_logic := '0';
  constant RTRTH_RSTVAL : std_logic_vector(3 downto 0) := x"0";
  constant ILBP_RSTVAL        : std_logic := '0';
  constant ENA_RSTVAL         : std_logic := '0';
  constant NISOFD_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- INT_STAT register
  --
  -- Reading this register returns logic 1 for each interrupt which was captured
  --  (interrupt vector). Writing logic 1 to any bit clears according bit of cap
  -- tured interrupt. Writing logic 0 has no effect.
  ------------------------------------------------------------------------------
  constant RXI_IND                : natural := 0;
  constant TXI_IND                : natural := 1;
  constant EWLI_IND               : natural := 2;
  constant DOI_IND                : natural := 3;
  constant EPI_IND                : natural := 4;
  constant ALI_IND                : natural := 5;
  constant BEI_IND                : natural := 6;
  constant LFI_IND                : natural := 7;
  constant RXFI_IND               : natural := 8;
  constant BSI_IND                : natural := 9;
  constant RBNEI_IND             : natural := 10;
  constant TXBHCI_IND            : natural := 11;

  -- INT_STAT register reset values
  constant RXI_RSTVAL         : std_logic := '0';
  constant TXI_RSTVAL         : std_logic := '0';
  constant EWLI_RSTVAL        : std_logic := '0';
  constant DOI_RSTVAL         : std_logic := '0';
  constant EPI_RSTVAL         : std_logic := '0';
  constant ALI_RSTVAL         : std_logic := '0';
  constant BEI_RSTVAL         : std_logic := '0';
  constant LFI_RSTVAL         : std_logic := '0';
  constant RXFI_RSTVAL        : std_logic := '0';
  constant BSI_RSTVAL         : std_logic := '0';
  constant RBNEI_RSTVAL       : std_logic := '0';
  constant TXBHCI_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- INT_ENA_SET register
  --
  -- Writing logic 1 to a bit enables according interrupt. Writing logic 0 has n
  -- o effect. Reading this register returns logic 1 for each enabled interrupt.
  --  If interrupt is captured in INT_STAT, enabled interrupt will cause "int" o
  -- utput to be asserted. Interrupts are level-based. To capture interrupt to I
  -- NT_STAT register, interrupt must be unmasked.
  ------------------------------------------------------------------------------
  constant INT_ENA_SET_L          : natural := 0;
  constant INT_ENA_SET_H         : natural := 11;

  -- INT_ENA_SET register reset values
  constant INT_ENA_SET_RSTVAL : std_logic_vector(11 downto 0) := x"000";

  ------------------------------------------------------------------------------
  -- INT_ENA_CLR register
  --
  -- Writing logic 1 disables according interrupt. Writing logic 0 has no effect
  -- . Reading this register has no effect. Disabled interrupt wil not affect "i
  -- nt" output of CAN Core event if it is captured in INT_STAT register.
  ------------------------------------------------------------------------------
  constant INT_ENA_CLR_L          : natural := 0;
  constant INT_ENA_CLR_H         : natural := 11;

  -- INT_ENA_CLR register reset values
  constant INT_ENA_CLR_RSTVAL : std_logic_vector(11 downto 0) := x"000";

  ------------------------------------------------------------------------------
  -- INT_MASK_SET register
  --
  -- Writing logic 1 masks according interrupt. Writing logic 0 has no effect. R
  -- eading this register returns logic 1 for each masked interrupt. If particul
  -- ar interrupt is masked, it won't be captured in INT_STAT register when inte
  -- rnal conditions for this interrupt are met (e.g RX Buffer is not empty for 
  -- RXNEI).
  ------------------------------------------------------------------------------
  constant INT_MASK_SET_L         : natural := 0;
  constant INT_MASK_SET_H        : natural := 11;

  -- INT_MASK_SET register reset values
  constant INT_MASK_SET_RSTVAL : std_logic_vector(11 downto 0) := x"000";

  ------------------------------------------------------------------------------
  -- INT_MASK_CLR register
  --
  -- Writing logic 1 un-masks according interrupt. Writing logic 0 has no effect
  -- . Reading this register has no effect. If particular interrupt is un-masked
  -- , it will be captured in INT_STAT register when internal conditions for thi
  -- s interrupt are met (e.g RX Buffer is not empty for RXNEI).
  ------------------------------------------------------------------------------
  constant INT_MASK_CLR_L         : natural := 0;
  constant INT_MASK_CLR_H        : natural := 11;

  -- INT_MASK_CLR register reset values
  constant INT_MASK_CLR_RSTVAL : std_logic_vector(11 downto 0) := x"000";

  ------------------------------------------------------------------------------
  -- BTR register
  --
  -- Bit timing register for nominal bit-rate. This register should be modified 
  -- only when SETTINGS[ENA]=0.
  ------------------------------------------------------------------------------
  constant PROP_L                 : natural := 0;
  constant PROP_H                 : natural := 6;
  constant PH1_L                  : natural := 7;
  constant PH1_H                 : natural := 12;
  constant PH2_L                 : natural := 13;
  constant PH2_H                 : natural := 18;
  constant BRP_L                 : natural := 19;
  constant BRP_H                 : natural := 26;
  constant SJW_L                 : natural := 27;
  constant SJW_H                 : natural := 31;

  -- BTR register reset values
  constant PROP_RSTVAL : std_logic_vector(6 downto 0) := "0000101";
  constant PH1_RSTVAL : std_logic_vector(5 downto 0) := "000011";
  constant PH2_RSTVAL : std_logic_vector(5 downto 0) := "000101";
  constant BRP_RSTVAL : std_logic_vector(7 downto 0) := x"0A";
  constant SJW_RSTVAL : std_logic_vector(4 downto 0) := "00010";

  ------------------------------------------------------------------------------
  -- BTR_FD register
  --
  -- Bit timing register for data bit-rate. This register should be modified onl
  -- y when SETTINGS[ENA]=0.
  ------------------------------------------------------------------------------
  constant PROP_FD_L              : natural := 0;
  constant PROP_FD_H              : natural := 5;
  constant PH1_FD_L               : natural := 7;
  constant PH1_FD_H              : natural := 11;
  constant PH2_FD_L              : natural := 13;
  constant PH2_FD_H              : natural := 17;
  constant BRP_FD_L              : natural := 19;
  constant BRP_FD_H              : natural := 26;
  constant SJW_FD_L              : natural := 27;
  constant SJW_FD_H              : natural := 31;

  -- BTR_FD register reset values
  constant PH2_FD_RSTVAL : std_logic_vector(4 downto 0) := "00011";
  constant PROP_FD_RSTVAL : std_logic_vector(5 downto 0) := "000011";
  constant PH1_FD_RSTVAL : std_logic_vector(4 downto 0) := "00011";
  constant BRP_FD_RSTVAL : std_logic_vector(7 downto 0) := x"04";
  constant SJW_FD_RSTVAL : std_logic_vector(4 downto 0) := "00010";

  ------------------------------------------------------------------------------
  -- EWL register
  --
  -- Error warning limit register. This register should be modified only when SE
  -- TTINGS[ENA]=0.
  ------------------------------------------------------------------------------
  constant EW_LIMIT_L             : natural := 0;
  constant EW_LIMIT_H             : natural := 7;

  -- EWL register reset values
  constant EW_LIMIT_RSTVAL : std_logic_vector(7 downto 0) := x"60";

  ------------------------------------------------------------------------------
  -- ERP register
  --
  -- Error passive limit register. This register should be modified only when SE
  -- TTINGS[ENA]=0.
  ------------------------------------------------------------------------------
  constant ERP_LIMIT_L            : natural := 8;
  constant ERP_LIMIT_H           : natural := 15;

  -- ERP register reset values
  constant ERP_LIMIT_RSTVAL : std_logic_vector(7 downto 0) := x"80";

  ------------------------------------------------------------------------------
  -- FAULT_STATE register
  --
  -- Fault confinement state of the node. This state can be manipulated by write
  -- s to CTR_PRES register. When these counters are set Fault confinement state
  --  changes automatically.
  ------------------------------------------------------------------------------
  constant ERA_IND               : natural := 16;
  constant ERP_IND               : natural := 17;
  constant BOF_IND               : natural := 18;

  -- FAULT_STATE register reset values
  constant ERP_RSTVAL         : std_logic := '0';
  constant BOF_RSTVAL         : std_logic := '0';
  constant ERA_RSTVAL         : std_logic := '1';

  ------------------------------------------------------------------------------
  -- RXC register
  --
  -- Counter for received frames.
  ------------------------------------------------------------------------------
  constant RXC_VAL_L              : natural := 0;
  constant RXC_VAL_H             : natural := 15;

  -- RXC register reset values
  constant RXC_VAL_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

  ------------------------------------------------------------------------------
  -- TXC register
  --
  -- Counter for transcieved frames.
  ------------------------------------------------------------------------------
  constant TXC_VAL_L             : natural := 16;
  constant TXC_VAL_H             : natural := 31;

  -- TXC register reset values
  constant TXC_VAL_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

  ------------------------------------------------------------------------------
  -- ERR_NORM register
  --
  ------------------------------------------------------------------------------
  constant ERR_NORM_VAL_L         : natural := 0;
  constant ERR_NORM_VAL_H        : natural := 15;

  -- ERR_NORM register reset values
  constant ERR_NORM_VAL_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

  ------------------------------------------------------------------------------
  -- ERR_FD register
  --
  ------------------------------------------------------------------------------
  constant ERR_FD_VAL_L          : natural := 16;
  constant ERR_FD_VAL_H          : natural := 31;

  -- ERR_FD register reset values
  constant ERR_FD_VAL_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

  ------------------------------------------------------------------------------
  -- CTR_PRES register
  --
  -- Register for manipulation with error counters.
  ------------------------------------------------------------------------------
  constant CTPV_L                 : natural := 0;
  constant CTPV_H                 : natural := 8;
  constant PTX_IND                : natural := 9;
  constant PRX_IND               : natural := 10;
  constant ENORM_IND             : natural := 11;
  constant EFD_IND               : natural := 12;

  -- CTR_PRES register reset values
  constant CTPV_RSTVAL : std_logic_vector(8 downto 0) := (OTHERS => '0');
  constant PTX_RSTVAL         : std_logic := '0';
  constant PRX_RSTVAL         : std_logic := '0';
  constant ENORM_RSTVAL       : std_logic := '0';
  constant EFD_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- FILTER_A_MASK register
  --
  -- Bit mask for acceptance filter A. The identifier format is the same as tran
  -- smitted and received identifier format. BASE Identifier is  in bits 28 : 18
  --  and Identifier extension are bits 17 : 0. Note that filter support is avai
  -- lable by default but it can be left out from synthesis (to save logic) by s
  -- etting "sup_filtA=false". If the particular filter is not supported, writes
  --  to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_MASK_A_VAL_L       : natural := 0;
  constant BIT_MASK_A_VAL_H      : natural := 28;

  -- FILTER_A_MASK register reset values
  constant BIT_MASK_A_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_A_VAL register
  --
  -- Bit value for acceptance filters. Filters A, B, C are available. The identi
  -- fier format is the same as transmitted and received identifier format. BASE
  --  Identifier is 11 LSB and Identifier extension are bits 28-12! Note that fi
  -- lter support is available by default but it can be left out from synthesis 
  -- (to save logic) by setting "sup_filtX=false";. If the particular filter is 
  -- not supported, writes to this register have no effect and read will return 
  -- all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_VAL_A_VAL_L        : natural := 0;
  constant BIT_VAL_A_VAL_H       : natural := 28;

  -- FILTER_A_VAL register reset values
  constant BIT_VAL_A_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_B_MASK register
  --
  -- Bit mask for acceptance filter B. The identifier format is the same as tran
  -- smitted and received identifier format. BASE Identifier is  in bits 28 : 18
  --  and Identifier extension are bits 17 : 0. Note that filter support is avai
  -- lable by default but it can be left out from synthesis (to save logic) by s
  -- etting "sup_filtB=false". If the particular filter is not supported, writes
  --  to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_MASK_B_VAL_L       : natural := 0;
  constant BIT_MASK_B_VAL_H      : natural := 28;

  -- FILTER_B_MASK register reset values
  constant BIT_MASK_B_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_B_VAL register
  --
  -- Bit value for acceptance filter B. The identifier format is the same as tra
  -- nsmitted and received identifier format. BASE Identifier is in bits 28 : 18
  --  and Identifier extension are bits 17 : 0. Note that filter support is avai
  -- lable by default but it can be left out from synthesis (to save logic) by s
  -- etting "sup_filtB=false". If the particular filter is not supported, writes
  --  to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_VAL_B_VAL_L        : natural := 0;
  constant BIT_VAL_B_VAL_H       : natural := 28;

  -- FILTER_B_VAL register reset values
  constant BIT_VAL_B_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_C_MASK register
  --
  -- Bit mask for acceptance filter C. The identifier format is the same as tran
  -- smitted and received identifier format. BASE Identifier is  in bits 28 : 18
  --  and Identifier extension are bits 17 : 0. Note that filter support is avai
  -- lable by default but it can be left out from synthesis (to save logic) by s
  -- etting "sup_filtC=false". If the particular filter is not supported, writes
  --  to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_MASK_C_VAL_L       : natural := 0;
  constant BIT_MASK_C_VAL_H      : natural := 28;

  -- FILTER_C_MASK register reset values
  constant BIT_MASK_C_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_C_VAL register
  --
  -- Bit value for acceptance filter C. The identifier format is the same as tra
  -- nsmitted and received identifier format. BASE Identifier is  in bits 28 : 1
  -- 8 and Identifier extension are bits 17 : 0. Note that filter support is ava
  -- ilable by default but it can be left out from synthesis (to save logic) by 
  -- setting "sup_filtC=false". If the particular filter is not supported, write
  -- s to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_VAL_C_VAL_L        : natural := 0;
  constant BIT_VAL_C_VAL_H       : natural := 28;

  -- FILTER_C_VAL register reset values
  constant BIT_VAL_C_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_RAN_LOW register
  --
  -- Low Identifier threshold for range filter. The identifier format is the sam
  -- e as transmitted and received identifier format. BASE Identifier is in bits
  --  28 : 18 and Identifier extension are bits 17 : 0. Note that filter support
  --  is available by default but it can be left out from synthesis (to save log
  -- ic) by setting "sup_range=false". If the particular filter is not supported
  -- , writes to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_RAN_LOW_VAL_L      : natural := 0;
  constant BIT_RAN_LOW_VAL_H     : natural := 28;

  -- FILTER_RAN_LOW register reset values
  constant BIT_RAN_LOW_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_RAN_HIGH register
  --
  -- High Identifier threshold for range filter. The identifier format is the sa
  -- me as transmitted and received identifier format. BASE Identifier is in bit
  -- s 28 : 18 and Identifier extension are bits 17 : 0. Note that filter suppor
  -- t is available by default but it can be left out from synthesis (to save lo
  -- gic) by setting "sup_range=false". If the particular filter is not supporte
  -- d, writes to this register have no effect and read will return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_RAN_HIGH_VAL_L     : natural := 0;
  constant BIT_RAN_HIGH_VAL_H    : natural := 28;

  -- FILTER_RAN_HIGH register reset values
  constant BIT_RAN_HIGH_VAL_RSTVAL
                 : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_CONTROL register
  --
  -- Every filter can be configured to accept only selected frame types. Every b
  -- it is active in logic 1.
  ------------------------------------------------------------------------------
  constant FANB_IND               : natural := 0;
  constant FANE_IND               : natural := 1;
  constant FAFB_IND               : natural := 2;
  constant FAFE_IND               : natural := 3;
  constant FBNB_IND               : natural := 4;
  constant FBNE_IND               : natural := 5;
  constant FBFB_IND               : natural := 6;
  constant FBFE_IND               : natural := 7;
  constant FCNB_IND               : natural := 8;
  constant FCNE_IND               : natural := 9;
  constant FCFB_IND              : natural := 10;
  constant FCFE_IND              : natural := 11;
  constant FRNB_IND              : natural := 12;
  constant FRNE_IND              : natural := 13;
  constant FRFB_IND              : natural := 14;
  constant FRFE_IND              : natural := 15;

  -- FILTER_CONTROL register reset values
  constant FANB_RSTVAL        : std_logic := '1';
  constant FAFB_RSTVAL        : std_logic := '1';
  constant FANE_RSTVAL        : std_logic := '1';
  constant FAFE_RSTVAL        : std_logic := '1';
  constant FBNB_RSTVAL        : std_logic := '0';
  constant FBNE_RSTVAL        : std_logic := '0';
  constant FBFB_RSTVAL        : std_logic := '0';
  constant FBFE_RSTVAL        : std_logic := '0';
  constant FCNB_RSTVAL        : std_logic := '0';
  constant FCNE_RSTVAL        : std_logic := '0';
  constant FCFB_RSTVAL        : std_logic := '0';
  constant FRFE_RSTVAL        : std_logic := '0';
  constant FRFB_RSTVAL        : std_logic := '0';
  constant FRNE_RSTVAL        : std_logic := '0';
  constant FRNB_RSTVAL        : std_logic := '0';
  constant FCFE_RSTVAL        : std_logic := '0';

  ------------------------------------------------------------------------------
  -- FILTER_STATUS register
  --
  -- This register provides information if the Core is synthesized with fillter 
  -- support.
  ------------------------------------------------------------------------------
  constant SFA_IND               : natural := 16;
  constant SFB_IND               : natural := 17;
  constant SFC_IND               : natural := 18;
  constant SFR_IND               : natural := 19;

  -- FILTER_STATUS register reset values

  ------------------------------------------------------------------------------
  -- RX_MEM_INFO register
  --
  -- Information register about FIFO memory of RX Buffer.
  ------------------------------------------------------------------------------
  constant RX_BUFF_SIZE_L         : natural := 0;
  constant RX_BUFF_SIZE_H        : natural := 12;
  constant RX_MEM_FREE_L         : natural := 16;
  constant RX_MEM_FREE_H         : natural := 28;

  -- RX_MEM_INFO register reset values

  ------------------------------------------------------------------------------
  -- RX_POINTERS register
  --
  -- Pointers in the RX FIFO buffer for read (by SW) and write (by Protocol cont
  -- rol FSM).
  ------------------------------------------------------------------------------
  constant RX_WPP_L               : natural := 0;
  constant RX_WPP_H              : natural := 11;
  constant RX_RPP_L              : natural := 16;
  constant RX_RPP_H              : natural := 27;

  -- RX_POINTERS register reset values
  constant RX_WPP_RSTVAL : std_logic_vector(11 downto 0) := x"000";
  constant RX_RPP_RSTVAL : std_logic_vector(11 downto 0) := x"000";

  ------------------------------------------------------------------------------
  -- RX_STATUS register
  --
  -- Information register one about FIFO Receive buffer.
  ------------------------------------------------------------------------------
  constant RXE_IND                : natural := 0;
  constant RXF_IND                : natural := 1;
  constant RXFRC_L                : natural := 4;
  constant RXFRC_H               : natural := 14;

  -- RX_STATUS register reset values
  constant RXE_RSTVAL         : std_logic := '1';
  constant RXF_RSTVAL         : std_logic := '1';
  constant RXFRC_RSTVAL : std_logic_vector(10 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_SETTINGS register
  --
  -- Settings register for FIFO RX Buffer.
  ------------------------------------------------------------------------------
  constant RTSOP_IND             : natural := 16;

  -- "RTSOP" field enumerated values
  constant RTS_END            : std_logic := '0';
  constant RTS_BEG            : std_logic := '1';

  -- RX_SETTINGS register reset values
  constant RTSOP_RSTVAL       : std_logic := '0';

  ------------------------------------------------------------------------------
  -- RX_DATA register
  --
  -- Read data word from RX Buffer.
  ------------------------------------------------------------------------------
  constant RX_DATA_L              : natural := 0;
  constant RX_DATA_H             : natural := 31;

  -- RX_DATA register reset values
  constant RX_DATA_RSTVAL : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- TX_STATUS register
  --
  -- Status of TXT Buffers. 
  ------------------------------------------------------------------------------
  constant TX1S_L                 : natural := 0;
  constant TX1S_H                 : natural := 3;
  constant TX2S_L                 : natural := 4;
  constant TX2S_H                 : natural := 7;
  constant TX3S_L                 : natural := 8;
  constant TX3S_H                : natural := 11;
  constant TX4S_L                : natural := 12;
  constant TX4S_H                : natural := 15;

  -- "TX1S" field enumerated values
  constant TXT_RDY : std_logic_vector(3 downto 0) := x"1";
  constant TXT_TRAN : std_logic_vector(3 downto 0) := x"2";
  constant TXT_ABTP : std_logic_vector(3 downto 0) := x"3";
  constant TXT_TOK : std_logic_vector(3 downto 0) := x"4";
  constant TXT_ERR : std_logic_vector(3 downto 0) := x"6";
  constant TXT_ABT : std_logic_vector(3 downto 0) := x"7";
  constant TXT_ETY : std_logic_vector(3 downto 0) := x"8";

  -- TX_STATUS register reset values
  constant TX2S_RSTVAL : std_logic_vector(3 downto 0) := x"8";
  constant TX1S_RSTVAL : std_logic_vector(3 downto 0) := x"8";
  constant TX3S_RSTVAL : std_logic_vector(3 downto 0) := x"8";
  constant TX4S_RSTVAL : std_logic_vector(3 downto 0) := x"8";

  ------------------------------------------------------------------------------
  -- TX_COMMAND register
  --
  -- Command register for TXT Buffers. Command is activated by setting TXC(E,R,A
  -- ) bit to logic 1. Buffer that receives the command is selected by setting b
  -- it TXBI(1..4) to logic 1. Command and index must be set by single access. R
  -- egister is automatically erased upon the command completion and 0 does not 
  -- need to be written. Reffer to description of TXT Buffer circuit for TXT buf
  -- fer State machine.   If TXCE and TXCR are applied simultaneously, only TXCE
  --  command is applied. If multiple commands are applied, only those which hav
  -- e effect in immediate state of the buffer are applied on a buffer.
  ------------------------------------------------------------------------------
  constant TXCE_IND               : natural := 0;
  constant TXCR_IND               : natural := 1;
  constant TXCA_IND               : natural := 2;
  constant TXB1_IND               : natural := 8;
  constant TXB2_IND               : natural := 9;
  constant TXB3_IND              : natural := 10;
  constant TXB4_IND              : natural := 11;

  -- TX_COMMAND register reset values
  constant TXCE_RSTVAL        : std_logic := '0';
  constant TXCR_RSTVAL        : std_logic := '0';
  constant TXCA_RSTVAL        : std_logic := '0';
  constant TXB1_RSTVAL        : std_logic := '0';
  constant TXB2_RSTVAL        : std_logic := '0';
  constant TXB3_RSTVAL        : std_logic := '0';
  constant TXB4_RSTVAL        : std_logic := '0';

  ------------------------------------------------------------------------------
  -- TX_PRIORITY register
  --
  -- Priority of the TXT Buffers in TX Arbitrator. Higher priority value signals
  --  that buffer is selected earlier for transmission. If two buffers have equa
  -- l priorities, the one with lower index is selected.
  ------------------------------------------------------------------------------
  constant TXT1P_L                : natural := 0;
  constant TXT1P_H                : natural := 2;
  constant TXT2P_L                : natural := 4;
  constant TXT2P_H                : natural := 6;
  constant TXT3P_L                : natural := 8;
  constant TXT3P_H               : natural := 10;
  constant TXT4P_L               : natural := 12;
  constant TXT4P_H               : natural := 14;

  -- TX_PRIORITY register reset values
  constant TXT1P_RSTVAL : std_logic_vector(2 downto 0) := "001";
  constant TXT2P_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant TXT3P_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant TXT4P_RSTVAL : std_logic_vector(2 downto 0) := "000";

  ------------------------------------------------------------------------------
  -- ERR_CAPT register
  --
  -- Last error frame capture.
  ------------------------------------------------------------------------------
  constant ERR_POS_L              : natural := 0;
  constant ERR_POS_H              : natural := 4;
  constant ERR_TYPE_L             : natural := 5;
  constant ERR_TYPE_H             : natural := 7;

  -- "ERR_POS" field enumerated values
  constant ERC_POS_SOF : std_logic_vector(4 downto 0) := "00000";
  constant ERC_POS_ARB : std_logic_vector(4 downto 0) := "00001";
  constant ERC_POS_CTRL : std_logic_vector(4 downto 0) := "00010";
  constant ERC_POS_DATA : std_logic_vector(4 downto 0) := "00011";
  constant ERC_POS_CRC : std_logic_vector(4 downto 0) := "00100";
  constant ERC_POS_ACK : std_logic_vector(4 downto 0) := "00101";
  constant ERC_POS_INTF : std_logic_vector(4 downto 0) := "00110";
  constant ERC_POS_ERR : std_logic_vector(4 downto 0) := "00111";
  constant ERC_POS_OVRL : std_logic_vector(4 downto 0) := "01000";
  constant ERC_POS_OTHER : std_logic_vector(4 downto 0) := "11111";

  -- "ERR_TYPE" field enumerated values
  constant ERC_BIT_ERR : std_logic_vector(2 downto 0) := "000";
  constant ERC_CRC_ERR : std_logic_vector(2 downto 0) := "001";
  constant ERC_FRM_ERR : std_logic_vector(2 downto 0) := "010";
  constant ERC_ACK_ERR : std_logic_vector(2 downto 0) := "011";
  constant ERC_STUF_ERR : std_logic_vector(2 downto 0) := "100";

  -- ERR_CAPT register reset values
  constant ERR_POS_RSTVAL : std_logic_vector(4 downto 0) := "11111";
  constant ERR_TYPE_RSTVAL : std_logic_vector(2 downto 0) := "000";

  ------------------------------------------------------------------------------
  -- ALC register
  --
  -- Arbitration lost capture register. Determines bit position of last arbitrat
  -- ion lost.
  ------------------------------------------------------------------------------
  constant ALC_BIT_L              : natural := 8;
  constant ALC_BIT_H             : natural := 12;
  constant ALC_ID_FIELD_L        : natural := 13;
  constant ALC_ID_FIELD_H        : natural := 15;

  -- "ALC_ID_FIELD" field enumerated values
  constant ALC_BASE_ID : std_logic_vector(2 downto 0) := "000";
  constant ALC_SRR_RTR : std_logic_vector(2 downto 0) := "001";
  constant ALC_IDE : std_logic_vector(2 downto 0) := "010";
  constant ALC_EXTENSION : std_logic_vector(2 downto 0) := "011";
  constant ALC_RTR : std_logic_vector(2 downto 0) := "100";

  -- ALC register reset values
  constant ALC_BIT_RSTVAL : std_logic_vector(4 downto 0) := "00000";
  constant ALC_ID_FIELD_RSTVAL : std_logic_vector(2 downto 0) := "000";

  ------------------------------------------------------------------------------
  -- TRV_DELAY register
  --
  ------------------------------------------------------------------------------
  constant TRV_DELAY_VALUE_L      : natural := 0;
  constant TRV_DELAY_VALUE_H     : natural := 15;

  -- TRV_DELAY register reset values
  constant TRV_DELAY_VALUE_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

  ------------------------------------------------------------------------------
  -- SSP_CFG register
  --
  -- Configuration of Secondary sampling point which is used for Transmitter in 
  -- Data Bit-Rate. This register should be modified only when SETTINGS[ENA]=0.
  ------------------------------------------------------------------------------
  constant SSP_OFFSET_L          : natural := 16;
  constant SSP_OFFSET_H          : natural := 22;
  constant SSP_SRC_L             : natural := 24;
  constant SSP_SRC_H             : natural := 25;

  -- "SSP_SRC" field enumerated values
  constant SSP_SRC_MEASURED : std_logic_vector(1 downto 0) := "00";
  constant SSP_SRC_MEAS_N_OFFSET : std_logic_vector(1 downto 0) := "01";
  constant SSP_SRC_OFFSET : std_logic_vector(1 downto 0) := "10";

  -- SSP_CFG register reset values
  constant SSP_OFFSET_RSTVAL : std_logic_vector(6 downto 0) := "0000000";
  constant SSP_SRC_RSTVAL : std_logic_vector(1 downto 0) := "00";

  ------------------------------------------------------------------------------
  -- RX_COUNTER register
  --
  -- Counter for received frames to enable bus traffic measurement
  ------------------------------------------------------------------------------
  constant RX_COUNTER_VAL_L       : natural := 0;
  constant RX_COUNTER_VAL_H      : natural := 31;

  -- RX_COUNTER register reset values
  constant RX_COUNTER_VAL_RSTVAL
                 : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- TX_COUNTER register
  --
  -- Counter for transmitted frames to enable bus traffic measurement.
  ------------------------------------------------------------------------------
  constant TX_COUNTER_VAL_L       : natural := 0;
  constant TX_COUNTER_VAL_H      : natural := 31;

  -- TX_COUNTER register reset values
  constant TX_COUNTER_VAL_RSTVAL
                 : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- DEBUG_REGISTER register
  --
  -- Register for reading out state of the controller. This register is only for
  --  debugging purposes!
  ------------------------------------------------------------------------------
  constant STUFF_COUNT_L          : natural := 0;
  constant STUFF_COUNT_H          : natural := 2;
  constant DESTUFF_COUNT_L        : natural := 3;
  constant DESTUFF_COUNT_H        : natural := 5;
  constant PC_ARB_IND             : natural := 6;
  constant PC_CON_IND             : natural := 7;
  constant PC_DAT_IND             : natural := 8;
  constant PC_CRC_IND             : natural := 9;
  constant PC_EOF_IND            : natural := 10;
  constant PC_OVR_IND            : natural := 11;
  constant PC_INT_IND            : natural := 12;

  -- DEBUG_REGISTER register reset values
  constant STUFF_COUNT_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant DESTUFF_COUNT_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant PC_ARB_RSTVAL      : std_logic := '0';
  constant PC_CON_RSTVAL      : std_logic := '0';
  constant PC_DAT_RSTVAL      : std_logic := '0';
  constant PC_CRC_RSTVAL      : std_logic := '0';
  constant PC_EOF_RSTVAL      : std_logic := '0';
  constant PC_OVR_RSTVAL      : std_logic := '0';
  constant PC_INT_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- YOLO_REG register
  --
  -- Register for fun :)
  ------------------------------------------------------------------------------
  constant YOLO_VAL_L             : natural := 0;
  constant YOLO_VAL_H            : natural := 31;

  -- YOLO_REG register reset values
  constant YOLO_VAL_RSTVAL : std_logic_vector(31 downto 0) := x"DEADBEEF";

  ------------------------------------------------------------------------------
  -- TIMESTAMP_LOW register
  --
  -- Register with mirrored values of timestamp input. Bits 31:0 of timestamp in
  -- put are available from this register. No synchronisation, nor shadowing is 
  -- implemented on TIMESTAMP_LOW/HIGH registers and user has to take care of pr
  -- oper read from both registers, since overflow of TIMESTAMP_LOW might occur 
  -- between read of TIMESTAMP_LOW and TIMESTAMP_HIGH.
  ------------------------------------------------------------------------------
  constant TIMESTAMP_LOW_L        : natural := 0;
  constant TIMESTAMP_LOW_H       : natural := 31;

  -- TIMESTAMP_LOW register reset values
  constant TIMESTAMP_LOW_RSTVAL : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- TIMESTAMP_HIGH register
  --
  -- Register with mirrored values of timestamp input. Bits 63:32 of timestamp i
  -- nput are available from this register. No synchronisation, nor shadowing is
  --  implemented on TIMESTAMP_LOW/HIGH registers and user has to take care of p
  -- roper read from both registers, since overflow of TIMESTAMP_LOW might occur
  --  between read of TIMESTAMP_LOW and TIMESTAMP_HIGH.
  ------------------------------------------------------------------------------
  constant TIMESTAMP_HIGH_L       : natural := 0;
  constant TIMESTAMP_HIGH_H      : natural := 31;

  -- TIMESTAMP_HIGH register reset values
  constant TIMESTAMP_HIGH_RSTVAL
                 : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- TXTB1_DATA_1 register
  --
  -- This adress word corresponds to FRAME_FORM word
  ------------------------------------------------------------------------------
  constant TXTB1_DATA_1_L         : natural := 0;
  constant TXTB1_DATA_1_H        : natural := 31;

  -- TXTB1_DATA_1 register reset values

  ------------------------------------------------------------------------------
  -- TXTB1_DATA_2 register
  --
  -- This adress word corresponds to IDENTIFIER word.
  ------------------------------------------------------------------------------
  constant TXTB1_DATA_2_L         : natural := 0;
  constant TXTB1_DATA_2_H        : natural := 31;

  -- TXTB1_DATA_2 register reset values

  ------------------------------------------------------------------------------
  -- TXTB1_DATA_20 register
  --
  -- This adress word corresponds to DATA_61_64 word.
  ------------------------------------------------------------------------------
  constant TXTB1_DATA_20_L        : natural := 0;
  constant TXTB1_DATA_20_H       : natural := 31;

  -- TXTB1_DATA_20 register reset values

  ------------------------------------------------------------------------------
  -- TXTB2_DATA_1 register
  --
  -- This adress word corresponds to FRAME_FORM word
  ------------------------------------------------------------------------------
  constant TXTB2_DATA_1_L         : natural := 0;
  constant TXTB2_DATA_1_H        : natural := 31;

  -- TXTB2_DATA_1 register reset values

  ------------------------------------------------------------------------------
  -- TXTB2_DATA_2 register
  --
  -- This adress word corresponds to IDENTIFIER word.
  ------------------------------------------------------------------------------
  constant TXTB2_DATA_2_L         : natural := 0;
  constant TXTB2_DATA_2_H        : natural := 31;

  -- TXTB2_DATA_2 register reset values

  ------------------------------------------------------------------------------
  -- TXTB2_DATA_20 register
  --
  -- This adress word corresponds to DATA_61_64 word.
  ------------------------------------------------------------------------------
  constant TXTB2_DATA_20_L        : natural := 0;
  constant TXTB2_DATA_20_H       : natural := 31;

  -- TXTB2_DATA_20 register reset values

  ------------------------------------------------------------------------------
  -- TXTB3_DATA_1 register
  --
  -- This adress word corresponds to FRAME_FORM word
  ------------------------------------------------------------------------------
  constant TXTB3_DATA_1_L         : natural := 0;
  constant TXTB3_DATA_1_H        : natural := 31;

  -- TXTB3_DATA_1 register reset values

  ------------------------------------------------------------------------------
  -- TXTB3_DATA_2 register
  --
  -- This adress word corresponds to IDENTIFIER word.
  ------------------------------------------------------------------------------
  constant TXTB3_DATA_2_L         : natural := 0;
  constant TXTB3_DATA_2_H        : natural := 31;

  -- TXTB3_DATA_2 register reset values

  ------------------------------------------------------------------------------
  -- TXTB3_DATA_20 register
  --
  -- This adress word corresponds to DATA_61_64 word.
  ------------------------------------------------------------------------------
  constant TXTB3_DATA_20_L        : natural := 0;
  constant TXTB3_DATA_20_H       : natural := 31;

  -- TXTB3_DATA_20 register reset values

  ------------------------------------------------------------------------------
  -- TXTB4_DATA_1 register
  --
  -- This adress word corresponds to FRAME_FORM word
  ------------------------------------------------------------------------------
  constant TXTB4_DATA_1_L         : natural := 0;
  constant TXTB4_DATA_1_H        : natural := 31;

  -- TXTB4_DATA_1 register reset values

  ------------------------------------------------------------------------------
  -- TXTB4_DATA_2 register
  --
  -- This adress word corresponds to IDENTIFIER word.
  ------------------------------------------------------------------------------
  constant TXTB4_DATA_2_L         : natural := 0;
  constant TXTB4_DATA_2_H        : natural := 31;

  -- TXTB4_DATA_2 register reset values

  ------------------------------------------------------------------------------
  -- TXTB4_DATA_20 register
  --
  -- This adress word corresponds to DATA_61_64 word.
  ------------------------------------------------------------------------------
  constant TXTB4_DATA_20_L        : natural := 0;
  constant TXTB4_DATA_20_H       : natural := 31;

  -- TXTB4_DATA_20 register reset values

  ------------------------------------------------------------------------------
  -- LOG_TRIG_CONFIG register
  --
  -- Register for configuration of event logging triggering conditions. If Event
  --  logger is in Ready state and any of triggering conditions appear it starts
  --  recording the events on the bus (moves to Running state). Logic 1 in each 
  -- bit means this triggering condition is valid.
  ------------------------------------------------------------------------------
  constant T_SOF_IND              : natural := 0;
  constant T_ARBL_IND             : natural := 1;
  constant T_REV_IND              : natural := 2;
  constant T_TRV_IND              : natural := 3;
  constant T_OVL_IND              : natural := 4;
  constant T_ERR_IND              : natural := 5;
  constant T_BRS_IND              : natural := 6;
  constant T_USRW_IND             : natural := 7;
  constant T_ARBS_IND             : natural := 8;
  constant T_CTRS_IND             : natural := 9;
  constant T_DATS_IND            : natural := 10;
  constant T_CRCS_IND            : natural := 11;
  constant T_ACKR_IND            : natural := 12;
  constant T_ACKNR_IND           : natural := 13;
  constant T_EWLR_IND            : natural := 14;
  constant T_ERPC_IND            : natural := 15;
  constant T_TRS_IND             : natural := 16;
  constant T_RES_IND             : natural := 17;

  -- LOG_TRIG_CONFIG register reset values
  constant T_SOF_RSTVAL       : std_logic := '0';
  constant T_ARBL_RSTVAL      : std_logic := '0';
  constant T_REV_RSTVAL       : std_logic := '0';
  constant T_TRV_RSTVAL       : std_logic := '0';
  constant T_OVL_RSTVAL       : std_logic := '0';
  constant T_RES_RSTVAL       : std_logic := '0';
  constant T_ERR_RSTVAL       : std_logic := '0';
  constant T_BRS_RSTVAL       : std_logic := '0';
  constant T_USRW_RSTVAL      : std_logic := '0';
  constant T_ARBS_RSTVAL      : std_logic := '0';
  constant T_CTRS_RSTVAL      : std_logic := '0';
  constant T_ACKNR_RSTVAL     : std_logic := '0';
  constant T_EWLR_RSTVAL      : std_logic := '0';
  constant T_ERPC_RSTVAL      : std_logic := '0';
  constant T_DATS_RSTVAL      : std_logic := '0';
  constant T_ACKR_RSTVAL      : std_logic := '0';
  constant T_TRS_RSTVAL       : std_logic := '0';
  constant T_CRCS_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_CAPT_CONFIG register
  --
  -- Register for configuring which events to capture by event logger into the l
  -- ogger FIFO memory when event logger is running.
  ------------------------------------------------------------------------------
  constant C_SOF_IND              : natural := 0;
  constant C_ARBL_IND             : natural := 1;
  constant C_REV_IND              : natural := 2;
  constant C_TRV_IND              : natural := 3;
  constant C_OVL_IND              : natural := 4;
  constant C_ERR_IND              : natural := 5;
  constant C_BRS_IND              : natural := 6;
  constant C_ARBS_IND             : natural := 7;
  constant C_CTRS_IND             : natural := 8;
  constant C_DATS_IND             : natural := 9;
  constant C_CRCS_IND            : natural := 10;
  constant C_ACKR_IND            : natural := 11;
  constant C_ACKNR_IND           : natural := 12;
  constant C_EWLR_IND            : natural := 13;
  constant C_ERC_IND             : natural := 14;
  constant C_TRS_IND             : natural := 15;
  constant C_RES_IND             : natural := 16;
  constant C_SYNE_IND            : natural := 17;
  constant C_STUFF_IND           : natural := 18;
  constant C_DESTUFF_IND         : natural := 19;
  constant C_OVR_IND             : natural := 20;

  -- LOG_CAPT_CONFIG register reset values
  constant C_SOF_RSTVAL       : std_logic := '0';
  constant C_ARBL_RSTVAL      : std_logic := '0';
  constant C_REV_RSTVAL       : std_logic := '0';
  constant C_TRV_RSTVAL       : std_logic := '0';
  constant C_OVL_RSTVAL       : std_logic := '0';
  constant C_ERR_RSTVAL       : std_logic := '0';
  constant C_BRS_RSTVAL       : std_logic := '0';
  constant C_ARBS_RSTVAL      : std_logic := '0';
  constant C_SYNE_RSTVAL      : std_logic := '0';
  constant C_STUFF_RSTVAL     : std_logic := '0';
  constant C_CTRS_RSTVAL      : std_logic := '0';
  constant C_DESTUFF_RSTVAL   : std_logic := '0';
  constant C_DATS_RSTVAL      : std_logic := '0';
  constant C_TRS_RSTVAL       : std_logic := '0';
  constant C_RES_RSTVAL       : std_logic := '0';
  constant C_OVR_RSTVAL       : std_logic := '0';
  constant C_CRCS_RSTVAL      : std_logic := '0';
  constant C_ACKR_RSTVAL      : std_logic := '0';
  constant C_ACKNR_RSTVAL     : std_logic := '0';
  constant C_EWLR_RSTVAL      : std_logic := '0';
  constant C_ERC_RSTVAL       : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_STATUS register
  --
  -- Status  register for Event logger.
  ------------------------------------------------------------------------------
  constant LOG_CFG_IND            : natural := 0;
  constant LOG_RDY_IND            : natural := 1;
  constant LOG_RUN_IND            : natural := 2;
  constant LOG_EXIST_IND          : natural := 7;
  constant LOG_SIZE_L             : natural := 8;
  constant LOG_SIZE_H            : natural := 15;

  -- LOG_STATUS register reset values
  constant LOG_CFG_RSTVAL     : std_logic := '1';
  constant LOG_RDY_RSTVAL     : std_logic := '0';
  constant LOG_RUN_RSTVAL     : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_POINTERS register
  --
  -- Pointers to Logger RAM memory.
  ------------------------------------------------------------------------------
  constant LOG_WPP_L             : natural := 16;
  constant LOG_WPP_H             : natural := 23;
  constant LOG_RPP_L             : natural := 24;
  constant LOG_RPP_H             : natural := 31;

  -- LOG_POINTERS register reset values
  constant LOG_WPP_RSTVAL : std_logic_vector(7 downto 0) := x"00";
  constant LOG_RPP_RSTVAL : std_logic_vector(7 downto 0) := x"00";

  ------------------------------------------------------------------------------
  -- LOG_COMMAND register
  --
  -- Register for controlling the state machine of Event logger and read pointer
  --  position. Every bit is active in logic 1.
  ------------------------------------------------------------------------------
  constant LOG_STR_IND            : natural := 0;
  constant LOG_ABT_IND            : natural := 1;
  constant LOG_UP_IND             : natural := 2;
  constant LOG_DOWN_IND           : natural := 3;

  -- LOG_COMMAND register reset values
  constant LOG_STR_RSTVAL     : std_logic := '0';
  constant LOG_ABT_RSTVAL     : std_logic := '0';
  constant LOG_UP_RSTVAL      : std_logic := '0';
  constant LOG_DOWN_RSTVAL    : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_CAPT_EVENT_1 register
  --
  -- First word of the captured event at read pointer position.
  ------------------------------------------------------------------------------
  constant EVENT_TS_48_16_L       : natural := 0;
  constant EVENT_TS_48_16_H      : natural := 31;

  -- LOG_CAPT_EVENT_1 register reset values
  constant EVENT_TS_48_16_RSTVAL
                 : std_logic_vector(31 downto 0) := x"00000000";

  ------------------------------------------------------------------------------
  -- LOG_CAPT_EVENT_2 register
  --
  -- Second word of the captured event at read pointer position.
  ------------------------------------------------------------------------------
  constant EVNT_TYPE_L            : natural := 0;
  constant EVNT_TYPE_H            : natural := 4;
  constant EVNT_DEN_L             : natural := 5;
  constant EVNT_DEN_H             : natural := 7;
  constant EVNT_DET_L             : natural := 8;
  constant EVNT_DET_H            : natural := 12;
  constant EVNT_DEA_L            : natural := 13;
  constant EVNT_DEA_H            : natural := 15;
  constant EVENT_TS_15_0_L       : natural := 16;
  constant EVENT_TS_15_0_H       : natural := 31;

  -- "EVNT_TYPE" field enumerated values
  constant SOF_EVNT : std_logic_vector(4 downto 0) := "00001";
  constant ARBL_EVNT : std_logic_vector(4 downto 0) := "00010";
  constant FREC_EVNT : std_logic_vector(4 downto 0) := "00011";
  constant TRANV_EVNT : std_logic_vector(4 downto 0) := "00100";
  constant OVRL_EVNT : std_logic_vector(4 downto 0) := "00101";
  constant ERR_EVNT : std_logic_vector(4 downto 0) := "00110";
  constant BRS_EVNT : std_logic_vector(4 downto 0) := "00111";
  constant ARBS_EVNT : std_logic_vector(4 downto 0) := "01000";
  constant CONS_EVNT : std_logic_vector(4 downto 0) := "01001";
  constant DATS_EVNT : std_logic_vector(4 downto 0) := "01010";
  constant CRCS_EVNT : std_logic_vector(4 downto 0) := "01011";
  constant ACKR_EVNT : std_logic_vector(4 downto 0) := "01100";
  constant ACKN_EVNT : std_logic_vector(4 downto 0) := "01101";
  constant EWLR_EVNT : std_logic_vector(4 downto 0) := "01110";
  constant FCSC_EVNT : std_logic_vector(4 downto 0) := "01111";
  constant TS_EVNT : std_logic_vector(4 downto 0) := "10000";
  constant RS_EVNT : std_logic_vector(4 downto 0) := "10001";
  constant SE_EVNT : std_logic_vector(4 downto 0) := "10010";
  constant STF_EVNT : std_logic_vector(4 downto 0) := "10011";
  constant DSTF_EVNT : std_logic_vector(4 downto 0) := "10100";
  constant DOR_EVNT : std_logic_vector(4 downto 0) := "10101";

  -- "EVNT_DET" field enumerated values
  constant ISN_FDSTF : std_logic_vector(4 downto 0) := "00000";
  constant ISN_FSTF : std_logic_vector(4 downto 0) := "00000";
  constant BIT_ERR : std_logic_vector(4 downto 0) := "00001";
  constant S_UP : std_logic_vector(4 downto 0) := "00001";
  constant IS_SYNC : std_logic_vector(4 downto 0) := "00001";
  constant IS_FDSTF : std_logic_vector(4 downto 0) := "00001";
  constant IS_FSTF : std_logic_vector(4 downto 0) := "00001";
  constant ST_ERR : std_logic_vector(4 downto 0) := "00010";
  constant S_DOWN : std_logic_vector(4 downto 0) := "00010";
  constant IS_PROP : std_logic_vector(4 downto 0) := "00010";
  constant CRC_ERR : std_logic_vector(4 downto 0) := "00100";
  constant IS_PH1 : std_logic_vector(4 downto 0) := "00100";
  constant ACK_ERR : std_logic_vector(4 downto 0) := "01000";
  constant IS_PH2 : std_logic_vector(4 downto 0) := "01000";
  constant FRM_ERR : std_logic_vector(4 downto 0) := "10000";

  -- "EVNT_DEA" field enumerated values
  constant NO_SNC : std_logic_vector(2 downto 0) := "000";
  constant HA_SNC : std_logic_vector(2 downto 0) := "001";
  constant RE_SNC : std_logic_vector(2 downto 0) := "010";

  -- LOG_CAPT_EVENT_2 register reset values
  constant EVNT_TYPE_RSTVAL : std_logic_vector(4 downto 0) := "00000";
  constant EVNT_DEN_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant EVNT_DET_RSTVAL : std_logic_vector(4 downto 0) := "00000";
  constant EVNT_DEA_RSTVAL : std_logic_vector(2 downto 0) := "000";
  constant EVENT_TS_15_0_RSTVAL : std_logic_vector(15 downto 0) := x"0000";

end package;
