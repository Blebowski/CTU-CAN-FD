--------------------------------------------------------------------------------
-- 
-- CAN with Flexible Data-Rate IP Core 
-- 
-- Copyright (C) 2017 Ondrej Ille <ondrej.ille@gmail.com>
-- 
-- Project advisor: Jiri Novak <jnovak@fel.cvut.cz>
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy 
-- of this VHDL component and associated documentation files (the "Component"), 
-- to deal in the Component without restriction, including without limitation 
-- the rights to use, copy, modify, merge, publish, distribute, sublicense, 
-- and/or sell copies of the Component, and to permit persons to whom the 
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in 
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE 
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER 
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS 
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents. 
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN 
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------
--------------------------------------------------------------------------------
-- Purpose:
-- Address constants for register map: CAN_FD_32bit_regsBit field constants fo
-- r register map: CAN_FD_8bit_regs. This file is autogenerated, do NOT edit!
--------------------------------------------------------------------------------

Library ieee;
use ieee.std_logic_1164.all;

package CAN_FD_register_map is

  ------------------------------------------------------------------------------
  -- DEVICE_ID register
  --
  -- The register contains an identifer of CAN FD IP function. It is used to det
  -- ermine whether CAN IP function is mapped correctly on its base address.
  ------------------------------------------------------------------------------
  constant DEVICE_ID_L            : natural := 0;
  constant DEVICE_ID_H           : natural := 31;

  --DEVICE_ID reset values
  constant DEVICE_ID_RSTVAL : std_logic_vector(31 downto 0) := x"0000cafd";

  ------------------------------------------------------------------------------
  -- MODE register
  --
  -- MODE register sets special operating modes of the controller. All bits are 
  -- active in logic 1.
  ------------------------------------------------------------------------------
  constant RST_IND                : natural := 0;
  constant STM_IND                : natural := 2;
  constant AFM_IND                : natural := 3;
  constant FDE_IND                : natural := 4;
  constant LOM_IND                : natural := 1;
  constant TSM_IND                : natural := 6;
  constant RTR_PREF_IND           : natural := 5;
  constant ACF_IND                : natural := 7;

  --MODE reset values
  constant RST_RSTVAL         : std_logic := '0';
  constant STM_RSTVAL         : std_logic := '0';
  constant AFM_RSTVAL         : std_logic := '0';
  constant FDE_RSTVAL         : std_logic := '1';
  constant LOM_RSTVAL         : std_logic := '0';
  constant TSM_RSTVAL         : std_logic := '0';
  constant RTR_PREF_RSTVAL    : std_logic := '1';
  constant ACF_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- COMMAND register
  --
  -- Writing logic 1 gives a command to the controller. The meaning of command i
  -- s different for every bit. This register is automatically erased when a com
  -- mand is finished.
  ------------------------------------------------------------------------------
  constant AT_IND                 : natural := 9;
  constant RRB_IND               : natural := 10;
  constant CDO_IND               : natural := 11;

  --COMMAND reset values
  constant AT_RSTVAL          : std_logic := '0';
  constant RRB_RSTVAL         : std_logic := '0';
  constant CDO_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- STATUS register
  --
  -- Register signals various states of CAN controller which are not mutually ex
  -- clusive. Every bit is active in logic 1.
  ------------------------------------------------------------------------------
  constant RBS_IND               : natural := 16;
  constant TBS_IND               : natural := 18;
  constant DOS_IND               : natural := 17;
  constant ET_IND                : natural := 19;
  constant RS_IND                : natural := 20;
  constant TS_IND                : natural := 21;
  constant ES_IND                : natural := 22;
  constant BS_IND                : natural := 23;

  --STATUS reset values
  constant RBS_RSTVAL         : std_logic := '0';
  constant TBS_RSTVAL         : std_logic := '0';
  constant DOS_RSTVAL         : std_logic := '0';
  constant ET_RSTVAL          : std_logic := '0';
  constant RS_RSTVAL          : std_logic := '0';
  constant TS_RSTVAL          : std_logic := '0';
  constant ES_RSTVAL          : std_logic := '0';
  constant BS_RSTVAL          : std_logic := '1';

  ------------------------------------------------------------------------------
  -- SETTINGS register
  --
  -- Register with enable bit of the controller.The configuration of retransmiss
  -- ion limit for failed frames is also located in this register. Furthermore c
  -- onfiguration of ISO FD CAN or CAN FD 1.0 is done here. Every bit is active 
  -- in logic 1.
  ------------------------------------------------------------------------------
  constant RTRLE_IND             : natural := 24;
  constant RTR_TH_L              : natural := 25;
  constant RTR_TH_H              : natural := 28;
  constant INT_LOOP_IND          : natural := 29;
  constant ENA_IND               : natural := 30;
  constant FD_TYPE_IND           : natural := 31;

  -- "ENA" field enumerated values
  constant DISABLED : std_logic := '0';
  constant ENABLED : std_logic := '1';

  -- "FD_TYPE" field enumerated values
  constant ISO_FD : std_logic := '0';
  constant NON_ISO_FD : std_logic := '1';

  --SETTINGS reset values
  constant RTRLE_RSTVAL       : std_logic := '0';
  constant RTR_TH_RSTVAL : std_logic_vector(3 downto 0) := (OTHERS => '0');
  constant INT_LOOP_RSTVAL    : std_logic := '0';
  constant ENA_RSTVAL         : std_logic := '0';
  constant FD_TYPE_RSTVAL     : std_logic := '0';

  ------------------------------------------------------------------------------
  -- INT register
  --
  -- This register contains interrupt vector of interrupts that were generated s
  -- ince the last read. If 8 bit or 16 bit access is executed to any of lowest 
  -- two bits the register is automatically erased.
  ------------------------------------------------------------------------------
  constant RI_IND                 : natural := 0;
  constant TI_IND                 : natural := 1;
  constant EI_IND                 : natural := 2;
  constant DOI_IND                : natural := 3;
  constant EPI_IND                : natural := 5;
  constant ALI_IND                : natural := 6;
  constant BEI_IND                : natural := 7;
  constant LFI_IND                : natural := 8;
  constant RFI_IND                : natural := 9;
  constant BSI_IND               : natural := 10;

  --INT reset values
  constant RI_RSTVAL          : std_logic := '0';
  constant TI_RSTVAL          : std_logic := '0';
  constant EI_RSTVAL          : std_logic := '0';
  constant DOI_RSTVAL         : std_logic := '0';
  constant EPI_RSTVAL         : std_logic := '0';
  constant ALI_RSTVAL         : std_logic := '0';
  constant BEI_RSTVAL         : std_logic := '0';
  constant LFI_RSTVAL         : std_logic := '0';
  constant RFI_RSTVAL         : std_logic := '0';
  constant BSI_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- INT_ENA register
  --
  -- Register enables interrupts by different sources. Logic 1 in each bit means
  --  interrupt is allowed
  ------------------------------------------------------------------------------
  constant EIE_IND               : natural := 18;
  constant DOIE_IND              : natural := 19;
  constant EPIE_IND              : natural := 21;
  constant ALIE_IND              : natural := 22;
  constant RIE_IND               : natural := 16;
  constant BEIE_IND              : natural := 23;
  constant LFIE_IND              : natural := 24;
  constant RFIE_IND              : natural := 25;
  constant BSIE_IND              : natural := 26;
  constant TIE_IND               : natural := 17;

  --INT_ENA reset values
  constant EIE_RSTVAL         : std_logic := '0';
  constant DOIE_RSTVAL        : std_logic := '0';
  constant EPIE_RSTVAL        : std_logic := '0';
  constant ALIE_RSTVAL        : std_logic := '0';
  constant RIE_RSTVAL         : std_logic := '0';
  constant BEIE_RSTVAL        : std_logic := '0';
  constant LFIE_RSTVAL        : std_logic := '0';
  constant RFIE_RSTVAL        : std_logic := '0';
  constant BSIE_RSTVAL        : std_logic := '0';
  constant TIE_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- BTR_FD register
  --
  -- Length of bit time segments for Data bit time in Time quanta. Note that SYN
  -- C segment always lasts one Time quanta.
  ------------------------------------------------------------------------------
  constant PH2_FD_L              : natural := 27;
  constant PH2_FD_H              : natural := 30;
  constant PROP_FD_L             : natural := 16;
  constant PROP_FD_H             : natural := 21;
  constant PH1_FD_L              : natural := 22;
  constant PH1_FD_H              : natural := 25;

  --BTR_FD reset values
  constant PH2_FD_RSTVAL : std_logic_vector(3 downto 0) := x"3";
  constant PROP_FD_RSTVAL : std_logic_vector(5 downto 0) := "000011";
  constant PH1_FD_RSTVAL : std_logic_vector(3 downto 0) := x"3";

  ------------------------------------------------------------------------------
  -- BTR register
  --
  -- The length of bit time segments for Nominal bit time in Time quanta. Note t
  -- hat SYNC segment always lasts one Time quanta.
  ------------------------------------------------------------------------------
  constant PROP_L                 : natural := 0;
  constant PROP_H                 : natural := 5;
  constant PH1_L                  : natural := 6;
  constant PH1_H                 : natural := 10;
  constant PH2_L                 : natural := 11;
  constant PH2_H                 : natural := 15;

  --BTR reset values
  constant PROP_RSTVAL : std_logic_vector(5 downto 0) := "000101";
  constant PH1_RSTVAL : std_logic_vector(4 downto 0) := "00011";
  constant PH2_RSTVAL : std_logic_vector(4 downto 0) := "00101";

  ------------------------------------------------------------------------------
  -- ALC register
  --
  -- Arbitration lost capture value
  ------------------------------------------------------------------------------
  constant ALC_VAL_L              : natural := 0;
  constant ALC_VAL_H              : natural := 4;

  --ALC reset values
  constant ALC_VAL_RSTVAL : std_logic_vector(4 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- SJW register
  --
  -- Synchronisation jump width registers for both Nominal and Data bit times.
  ------------------------------------------------------------------------------
  constant SJW_L                  : natural := 8;
  constant SJW_H                 : natural := 11;
  constant SJW_FD_L              : natural := 12;
  constant SJW_FD_H              : natural := 15;

  --SJW reset values
  constant SJW_RSTVAL : std_logic_vector(3 downto 0) := x"2";
  constant SJW_FD_RSTVAL : std_logic_vector(3 downto 0) := x"2";

  ------------------------------------------------------------------------------
  -- BRP register
  --
  -- Baud rate Prescaler register for Nominal bit time. Specifies time quanta du
  -- ration.
  ------------------------------------------------------------------------------
  constant BRP_L                 : natural := 16;
  constant BRP_H                 : natural := 21;

  --BRP reset values
  constant BRP_RSTVAL : std_logic_vector(5 downto 0) := "001010";

  ------------------------------------------------------------------------------
  -- BRP_FD register
  --
  -- Baud rate Prescaler register for Data bit time. Specifies time quanta durat
  -- ion.
  ------------------------------------------------------------------------------
  constant BRP_FD_L              : natural := 24;
  constant BRP_FD_H              : natural := 29;

  --BRP_FD reset values
  constant BRP_FD_RSTVAL : std_logic_vector(5 downto 0) := "000100";

  ------------------------------------------------------------------------------
  -- EWL register
  --
  -- Error warning limit register. If an error warning limit is reached interrup
  -- t can be called. Error warning limit indicatea heavily disturbed bus. Note 
  -- that according to CAN specification this value is fixed at 96 and should no
  -- t be configurable! The configuration of this value is one of the extra feat
  -- ures of this IP Core.
  ------------------------------------------------------------------------------
  constant EWL_LIMIT_L            : natural := 0;
  constant EWL_LIMIT_H            : natural := 7;

  --EWL reset values
  constant EWL_LIMIT_RSTVAL : std_logic_vector(7 downto 0) := x"60";

  ------------------------------------------------------------------------------
  -- ERP register
  --
  -- Error passive limit. When one of error counters (RXC/TXC) exceeds this valu
  -- e, it changes Fault confinement state to error passive. Note that according
  --  to CAN specification this value is fixed at 128 and should not be configur
  -- able! The configuration of this value is one of the extra features of this 
  -- IP Core. Note that IP Core always turns to bus_off state once any error cou
  -- nter reaches 255!
  ------------------------------------------------------------------------------
  constant ERP_LIMIT_L            : natural := 8;
  constant ERP_LIMIT_H           : natural := 15;

  --ERP reset values
  constant ERP_LIMIT_RSTVAL : std_logic_vector(7 downto 0) := x"80";

  ------------------------------------------------------------------------------
  -- FAULT_STATE register
  --
  -- Fault confinement state of the node. This state can be manipulated by writi
  -- ng into registers RXC/TXC and ERP_LIMIT of ERP register. When these counter
  -- s are set Fault confinement state changes automatically.
  ------------------------------------------------------------------------------
  constant ERP_IND               : natural := 17;
  constant BOF_IND               : natural := 18;
  constant ERA_IND               : natural := 16;

  --FAULT_STATE reset values
  constant ERP_RSTVAL         : std_logic := '0';
  constant BOF_RSTVAL         : std_logic := '0';
  constant ERA_RSTVAL         : std_logic := '1';

  ------------------------------------------------------------------------------
  -- FILTER_A_VAL register
  --
  -- Bit value for acceptance filters. Filters A, B, C are available. The identi
  -- fier format is the same as transmitted and received identifier format. BASE
  --  Identifier is 11 LSB and Identifier extension are bits 28-12! Note that fi
  -- lter support is available by default but it can be left out from synthesis 
  -- (to save logic) by setting "sup_filtX=false";. If the particular filter is 
  -- not supported, writes to this register have no effect and read will return 
  -- all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_VAL_A_VAL_L        : natural := 0;
  constant BIT_VAL_A_VAL_H       : natural := 28;

  --FILTER_A_VAL reset values
  constant BIT_VAL_A_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_STATUS register
  --
  -- This register provides information about whether the Core is synthesized wi
  -- th fillter support.
  ------------------------------------------------------------------------------
  constant SUP_FILTA_IND         : natural := 16;
  constant SUP_FILTB_IND         : natural := 17;
  constant SUP_RANGE_IND         : natural := 19;
  constant SUP_FILTC_IND         : natural := 18;

  --FILTER_STATUS reset values

  ------------------------------------------------------------------------------
  -- RX_MF register
  --
  -- Number of free (32 bit) words in RX Buffer
  ------------------------------------------------------------------------------
  constant RX_MF_VALUE_L         : natural := 16;
  constant RX_MF_VALUE_H         : natural := 23;

  --RX_MF reset values

  ------------------------------------------------------------------------------
  -- RX_MC register
  --
  -- Register with number of frames in the receive buffer.
  ------------------------------------------------------------------------------
  constant RX_MC_VALUE_L          : natural := 8;
  constant RX_MC_VALUE_H         : natural := 15;

  --RX_MC reset values

  ------------------------------------------------------------------------------
  -- TX_SETTINGS register
  --
  -- This register controls the access into TX buffers. All bits are active in l
  -- ogic 1.
  ------------------------------------------------------------------------------
  constant TXT1_ALLOW_IND         : natural := 0;
  constant TXT2_ALLOW_IND         : natural := 1;
  constant BUF_DIR_IND            : natural := 2;
  constant FRAME_SWAP_IND         : natural := 3;

  --TX_SETTINGS reset values
  constant TXT1_ALLOW_RSTVAL  : std_logic := '1';
  constant TXT2_ALLOW_RSTVAL  : std_logic := '1';
  constant BUF_DIR_RSTVAL     : std_logic := '0';
  constant FRAME_SWAP_RSTVAL  : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_TRIG_CONFIG register
  --
  -- Register for configuration of event logging triggering conditions. If Event
  --  logger is in Ready state and any of triggering conditions appear it starts
  --  recording the events on the bus (moves to Running state). Logic 1 in each 
  -- bit means this triggering condition is valid.
  ------------------------------------------------------------------------------
  constant T_SOF_IND              : natural := 0;
  constant T_ARBL_IND             : natural := 1;
  constant T_TRV_IND              : natural := 3;
  constant T_REV_IND              : natural := 2;
  constant T_ERPC_IND            : natural := 15;
  constant T_OVL_IND              : natural := 4;
  constant T_ERR_IND              : natural := 5;
  constant T_BRS_IND              : natural := 6;
  constant T_TRS_IND             : natural := 16;
  constant T_USRW_IND             : natural := 7;
  constant T_EWLR_IND            : natural := 14;
  constant T_ARBS_IND             : natural := 8;
  constant T_CTRS_IND             : natural := 9;
  constant T_ACKNR_IND           : natural := 13;
  constant T_RES_IND             : natural := 17;
  constant T_ACKR_IND            : natural := 12;
  constant T_DATS_IND            : natural := 10;
  constant T_CRCS_IND            : natural := 11;

  --LOG_TRIG_CONFIG reset values
  constant T_SOF_RSTVAL       : std_logic := '0';
  constant T_ARBL_RSTVAL      : std_logic := '0';
  constant T_TRV_RSTVAL       : std_logic := '0';
  constant T_REV_RSTVAL       : std_logic := '0';
  constant T_ERPC_RSTVAL      : std_logic := '0';
  constant T_OVL_RSTVAL       : std_logic := '0';
  constant T_ERR_RSTVAL       : std_logic := '0';
  constant T_BRS_RSTVAL       : std_logic := '0';
  constant T_TRS_RSTVAL       : std_logic := '0';
  constant T_USRW_RSTVAL      : std_logic := '0';
  constant T_EWLR_RSTVAL      : std_logic := '0';
  constant T_ARBS_RSTVAL      : std_logic := '0';
  constant T_CTRS_RSTVAL      : std_logic := '0';
  constant T_ACKNR_RSTVAL     : std_logic := '0';
  constant T_RES_RSTVAL       : std_logic := '0';
  constant T_ACKR_RSTVAL      : std_logic := '0';
  constant T_DATS_RSTVAL      : std_logic := '0';
  constant T_CRCS_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_WPP register
  --
  ------------------------------------------------------------------------------
  constant LOG_WPP_VAL_L         : natural := 16;
  constant LOG_WPP_VAL_H         : natural := 23;

  --LOG_WPP reset values
  constant LOG_WPP_VAL_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- LOG_STATUS register
  --
  -- Status  register for Event logger.
  ------------------------------------------------------------------------------
  constant LOG_CFG_IND            : natural := 0;
  constant LOG_RDY_IND            : natural := 1;
  constant LOG_RUN_IND            : natural := 2;
  constant LOG_EXIST_IND          : natural := 7;
  constant LOG_SIZE_L             : natural := 8;
  constant LOG_SIZE_H            : natural := 15;

  --LOG_STATUS reset values
  constant LOG_CFG_RSTVAL     : std_logic := '1';
  constant LOG_RDY_RSTVAL     : std_logic := '0';
  constant LOG_RUN_RSTVAL     : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_CAPT_EVENT_2 register
  --
  -- Second word of the logged event details.
  ------------------------------------------------------------------------------
  constant EVENT_TS_15_0_L       : natural := 16;
  constant EVENT_TS_15_0_H       : natural := 31;
  constant EVENT_DETAILS_L        : natural := 8;
  constant EVENT_DETAILS_H       : natural := 15;
  constant EVENT_TYPE_L           : natural := 0;
  constant EVENT_TYPE_H           : natural := 7;

  -- "EVENT_TYPE" field enumerated values
  constant SOF_EVNT : std_logic_vector(7 downto 0) := "00000001";
  constant ALO_EVNT : std_logic_vector(7 downto 0) := "00000010";
  constant REC_EVNT : std_logic_vector(7 downto 0) := "00000011";
  constant TRAN_EVNT : std_logic_vector(7 downto 0) := "00000100";
  constant OVLD_EVNT : std_logic_vector(7 downto 0) := "00000101";
  constant ERR_EVNT : std_logic_vector(7 downto 0) := "00000110";
  constant BRS_EVNT : std_logic_vector(7 downto 0) := "00000111";
  constant ARB_EVNT : std_logic_vector(7 downto 0) := "00001000";
  constant CTRL_EVNT : std_logic_vector(7 downto 0) := "00001001";
  constant DATA_EVNT : std_logic_vector(7 downto 0) := "00001010";
  constant CRC_EVNT : std_logic_vector(7 downto 0) := "00001011";
  constant ACK_EVNT : std_logic_vector(7 downto 0) := "00001100";
  constant NACK_EVNT : std_logic_vector(7 downto 0) := "00001101";
  constant EWL_EVNT : std_logic_vector(7 downto 0) := "00001110";
  constant ERP_EVNT : std_logic_vector(7 downto 0) := "00001111";
  constant TXS_EVNT : std_logic_vector(7 downto 0) := "00010000";
  constant RXS_EVNT : std_logic_vector(7 downto 0) := "00010001";
  constant SYNC_EVNT : std_logic_vector(7 downto 0) := "00010010";
  constant STUF_EVNT : std_logic_vector(7 downto 0) := "00010011";
  constant DSTF_EVNT : std_logic_vector(7 downto 0) := "00010100";
  constant OVR_EVNT : std_logic_vector(7 downto 0) := "00010101";

  --LOG_CAPT_EVENT_2 reset values
  constant EVENT_TS_15_0_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');
  constant EVENT_DETAILS_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');
  constant EVENT_TYPE_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- LOG_CAPT_EVENT_1 register
  --
  -- First word of the logged event details.
  ------------------------------------------------------------------------------
  constant EVENT_TIME_STAMP_47_TO_16_L : natural := 0;
  constant EVENT_TIME_STAMP_47_TO_16_H : natural := 31;

  --LOG_CAPT_EVENT_1 reset values
  constant EVENT_TIME_STAMP_47_TO_16_RSTVAL : std_logic_vector(31 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- YOLO_REG register
  --
  -- Register for fun :)
  ------------------------------------------------------------------------------
  constant YOLO_VAL_L             : natural := 0;
  constant YOLO_VAL_H            : natural := 31;

  --YOLO_REG reset values
  constant YOLO_VAL_RSTVAL : std_logic_vector(31 downto 0) := x"deadbeef";

  ------------------------------------------------------------------------------
  -- DEBUG_REGISTER register
  --
  -- Register for reading out state of the controller. This register is only for
  --  debugging purposes!
  ------------------------------------------------------------------------------
  constant STUFF_COUNT_L          : natural := 0;
  constant STUFF_COUNT_H          : natural := 2;
  constant DESTUFF_COUNT_L        : natural := 3;
  constant DESTUFF_COUNT_H        : natural := 5;
  constant PC_ARB_IND             : natural := 6;
  constant PC_CON_IND             : natural := 7;
  constant PC_DAT_IND             : natural := 8;
  constant PC_CRC_IND             : natural := 9;
  constant PC_EOF_IND            : natural := 10;
  constant PC_OVR_IND            : natural := 11;
  constant PC_INT_IND            : natural := 12;

  --DEBUG_REGISTER reset values
  constant STUFF_COUNT_RSTVAL : std_logic_vector(2 downto 0) := (OTHERS => '0');
  constant DESTUFF_COUNT_RSTVAL : std_logic_vector(2 downto 0) := (OTHERS => '0');
  constant PC_ARB_RSTVAL      : std_logic := '0';
  constant PC_CON_RSTVAL      : std_logic := '0';
  constant PC_DAT_RSTVAL      : std_logic := '0';
  constant PC_CRC_RSTVAL      : std_logic := '0';
  constant PC_EOF_RSTVAL      : std_logic := '0';
  constant PC_OVR_RSTVAL      : std_logic := '0';
  constant PC_INT_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_COMMAND register
  --
  -- Register for controlling the state machine of Event logger and read pointer
  --  position. Every bit is active in logic 1.
  ------------------------------------------------------------------------------
  constant LOG_STR_IND            : natural := 0;
  constant LOG_ABT_IND            : natural := 1;
  constant LOG_UP_IND             : natural := 2;
  constant LOG_DOWN_IND           : natural := 3;

  --LOG_COMMAND reset values
  constant LOG_STR_RSTVAL     : std_logic := '0';
  constant LOG_ABT_RSTVAL     : std_logic := '0';
  constant LOG_UP_RSTVAL      : std_logic := '0';
  constant LOG_DOWN_RSTVAL    : std_logic := '0';

  ------------------------------------------------------------------------------
  -- LOG_RPP register
  --
  ------------------------------------------------------------------------------
  constant LOG_RPP_VAL_L         : natural := 24;
  constant LOG_RPP_VAL_H         : natural := 31;

  --LOG_RPP reset values
  constant LOG_RPP_VAL_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- LOG_CAPT_CONFIG register
  --
  -- Register for configuring which events to capture by event logger into the l
  -- ogger FIFO memory when event logger is running.
  ------------------------------------------------------------------------------
  constant C_SOF_IND              : natural := 0;
  constant C_ARBL_IND             : natural := 1;
  constant C_REV_IND              : natural := 2;
  constant C_TRV_IND              : natural := 3;
  constant C_OVL_IND              : natural := 4;
  constant C_DESTUFF_IND         : natural := 19;
  constant C_ERR_IND              : natural := 5;
  constant C_BRS_IND              : natural := 6;
  constant C_STUFF_IND           : natural := 18;
  constant C_SYNE_IND            : natural := 17;
  constant C_RES_IND             : natural := 16;
  constant C_ACKNR_IND           : natural := 12;
  constant C_OVR_IND             : natural := 20;
  constant C_EWLR_IND            : natural := 13;
  constant C_ARBS_IND             : natural := 7;
  constant C_CTRS_IND             : natural := 8;
  constant C_ERC_IND             : natural := 14;
  constant C_DATS_IND             : natural := 9;
  constant C_ACKR_IND            : natural := 11;
  constant C_TRS_IND             : natural := 15;
  constant C_CRCS_IND            : natural := 10;

  --LOG_CAPT_CONFIG reset values
  constant C_SOF_RSTVAL       : std_logic := '0';
  constant C_ARBL_RSTVAL      : std_logic := '0';
  constant C_REV_RSTVAL       : std_logic := '0';
  constant C_TRV_RSTVAL       : std_logic := '0';
  constant C_OVL_RSTVAL       : std_logic := '0';
  constant C_DESTUFF_RSTVAL   : std_logic := '0';
  constant C_ERR_RSTVAL       : std_logic := '0';
  constant C_BRS_RSTVAL       : std_logic := '0';
  constant C_STUFF_RSTVAL     : std_logic := '0';
  constant C_SYNE_RSTVAL      : std_logic := '0';
  constant C_RES_RSTVAL       : std_logic := '0';
  constant C_ACKNR_RSTVAL     : std_logic := '0';
  constant C_OVR_RSTVAL       : std_logic := '0';
  constant C_EWLR_RSTVAL      : std_logic := '0';
  constant C_ARBS_RSTVAL      : std_logic := '0';
  constant C_CTRS_RSTVAL      : std_logic := '0';
  constant C_ERC_RSTVAL       : std_logic := '0';
  constant C_DATS_RSTVAL      : std_logic := '0';
  constant C_ACKR_RSTVAL      : std_logic := '0';
  constant C_TRS_RSTVAL       : std_logic := '0';
  constant C_CRCS_RSTVAL      : std_logic := '0';

  ------------------------------------------------------------------------------
  -- TX_COUNTER register
  --
  -- Counter for transmitted frames to enable bus traffic measurement
  ------------------------------------------------------------------------------
  constant TX_COUNTER_VAL_L       : natural := 0;
  constant TX_COUNTER_VAL_H      : natural := 31;

  --TX_COUNTER reset values
  constant TX_COUNTER_VAL_RSTVAL : std_logic_vector(31 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_COUNTER register
  --
  -- Counter for received frames to enable bus traffic measurement
  ------------------------------------------------------------------------------
  constant RX_COUNTER_VAL_L       : natural := 0;
  constant RX_COUNTER_VAL_H      : natural := 31;

  --RX_COUNTER reset values
  constant RX_COUNTER_VAL_RSTVAL : std_logic_vector(31 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- ERR_CAPT register
  --
  -- Last error frame capture.
  ------------------------------------------------------------------------------
  constant ERR_POS_L              : natural := 0;
  constant ERR_POS_H              : natural := 4;
  constant ERR_TYPE_L             : natural := 5;
  constant ERR_TYPE_H             : natural := 7;

  -- "ERR_POS" field enumerated values
  constant ERC_POS_SOF : std_logic_vector(4 downto 0) := "00000";
  constant ERC_POS_ARB : std_logic_vector(4 downto 0) := "00001";
  constant ERC_POS_CTRL : std_logic_vector(4 downto 0) := "00010";
  constant ERC_POS_DATA : std_logic_vector(4 downto 0) := "00011";
  constant ERC_POS_CRC : std_logic_vector(4 downto 0) := "00100";
  constant ERC_POS_ACK : std_logic_vector(4 downto 0) := "00101";
  constant ERC_POS_INTF : std_logic_vector(4 downto 0) := "00110";
  constant ERC_POS_ERR : std_logic_vector(4 downto 0) := "00111";
  constant ERC_POS_OVRL : std_logic_vector(4 downto 0) := "01000";
  constant ERC_POS_OTHER : std_logic_vector(4 downto 0) := "11111";

  -- "ERR_TYPE" field enumerated values
  constant ERC_BIT_ERR : std_logic_vector(2 downto 0) := "000";
  constant ERC_CRC_ERR : std_logic_vector(2 downto 0) := "001";
  constant ERC_FRM_ERR : std_logic_vector(2 downto 0) := "010";
  constant ERC_ACK_ERR : std_logic_vector(2 downto 0) := "011";
  constant ERC_STUF_ERR : std_logic_vector(2 downto 0) := "100";

  --ERR_CAPT reset values
  constant ERR_POS_RSTVAL : std_logic_vector(4 downto 0) := "11111";
  constant ERR_TYPE_RSTVAL : std_logic_vector(2 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- TX_STATUS register
  --
  -- Status of the TXT Buffers
  ------------------------------------------------------------------------------
  constant TXT2_EMPTY_IND         : natural := 1;
  constant TXT1_EMPTY_IND         : natural := 0;
  constant TX_TIME_SUPPORT_IND    : natural := 2;

  --TX_STATUS reset values
  constant TXT2_EMPTY_RSTVAL  : std_logic := '1';
  constant TXT1_EMPTY_RSTVAL  : std_logic := '1';

  ------------------------------------------------------------------------------
  -- TRV_DELAY register
  --
  ------------------------------------------------------------------------------
  constant TRV_DELAY_VALUE_L      : natural := 0;
  constant TRV_DELAY_VALUE_H     : natural := 15;

  --TRV_DELAY reset values
  constant TRV_DELAY_VALUE_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_DATA register
  --
  -- The recieve buffer data at read pointer position in FIFO. CAN Frame layout 
  -- in RX buffer is described in Figure 7. By reading data from this register r
  -- ead_pointer is automatically increased, as long as there is next data word 
  -- stored in the buffer. Next Read from this register returns next word of CAN
  --  frame. First stored word in the buffer is FRAME_FORM, next TIMESTAMP_U etc
  -- . In detail bits of each word have following meaning. If any access is exec
  -- uted (8 bit, 16 bit or 32 bit), the read_pointer automatically increases. I
  -- t is recomended to use 32 bit acccess on this register.
  ------------------------------------------------------------------------------
  constant RX_DATA_L              : natural := 0;
  constant RX_DATA_H             : natural := 31;

  --RX_DATA reset values
  constant RX_DATA_RSTVAL : std_logic_vector(31 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_RPP register
  --
  -- Read pointer position in th Receive buffer. When a new frame is stored writ
  -- e pointer is increased accordingly.
  ------------------------------------------------------------------------------
  constant RX_RPP_VAL_L          : natural := 16;
  constant RX_RPP_VAL_H          : natural := 23;

  --RX_RPP reset values
  constant RX_RPP_VAL_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_WPP register
  --
  -- Write pointer position in th Receive buffer. When a new frame is stored wri
  -- te pointer is increased
  ------------------------------------------------------------------------------
  constant RX_WPP_VALUE_L         : natural := 8;
  constant RX_WPP_VALUE_H        : natural := 15;

  --RX_WPP reset values
  constant RX_WPP_VALUE_RSTVAL : std_logic_vector(7 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RX_BUFF_SIZE register
  --
  -- Size of th Receive buffer. This parameter is configurable before synthesis.
  ------------------------------------------------------------------------------
  constant RX_BUFF_SIZE_VALUE_L   : natural := 0;
  constant RX_BUFF_SIZE_VALUE_H   : natural := 7;

  --RX_BUFF_SIZE reset values

  ------------------------------------------------------------------------------
  -- RX_STATUS register
  --
  -- Information register one about FIFO Receive buffer.
  ------------------------------------------------------------------------------
  constant RX_EMPTY_IND           : natural := 0;
  constant RX_FULL_IND            : natural := 1;

  --RX_STATUS reset values
  constant RX_EMPTY_RSTVAL    : std_logic := '1';
  constant RX_FULL_RSTVAL     : std_logic := '1';

  ------------------------------------------------------------------------------
  -- FILTER_CONTROL register
  --
  -- Every filter can be set to accept only selected frame types. Every bit acti
  -- ve in logic 1.
  ------------------------------------------------------------------------------
  constant FILT_A_BASIC_IND       : natural := 0;
  constant FILT_A_FD_BAS_IND      : natural := 2;
  constant FILT_A_EXT_IND         : natural := 1;
  constant FILT_A_FD_EXT_IND      : natural := 3;
  constant FILT_B_BASIC_IND       : natural := 4;
  constant FILT_B_EXT_IND         : natural := 5;
  constant FILT_B_FD_BAS_IND      : natural := 6;
  constant FILT_B_FD_EXT_IND      : natural := 7;
  constant FILT_C_BASIC_IND       : natural := 8;
  constant FILT_C_EXT_IND         : natural := 9;
  constant FILT_C_FD_BAS_IND     : natural := 10;
  constant FILT_RANGE_FD_EXT_IND : natural := 15;
  constant FILT_RANGE_FD_BAS_IND : natural := 14;
  constant FILT_RANGE_EXT_IND    : natural := 13;
  constant FILT_RANGE_BASIC_IND  : natural := 12;
  constant FILT_C_FD_EXT_IND     : natural := 11;

  --FILTER_CONTROL reset values
  constant FILT_A_BASIC_RSTVAL : std_logic := '1';
  constant FILT_A_FD_BAS_RSTVAL : std_logic := '1';
  constant FILT_A_EXT_RSTVAL  : std_logic := '1';
  constant FILT_A_FD_EXT_RSTVAL : std_logic := '1';
  constant FILT_B_BASIC_RSTVAL : std_logic := '0';
  constant FILT_B_EXT_RSTVAL  : std_logic := '0';
  constant FILT_B_FD_BAS_RSTVAL : std_logic := '0';
  constant FILT_B_FD_EXT_RSTVAL : std_logic := '0';
  constant FILT_C_BASIC_RSTVAL : std_logic := '0';
  constant FILT_C_EXT_RSTVAL  : std_logic := '0';
  constant FILT_C_FD_BAS_RSTVAL : std_logic := '0';
  constant FILT_RANGE_FD_EXT_RSTVAL : std_logic := '0';
  constant FILT_RANGE_FD_BAS_RSTVAL : std_logic := '0';
  constant FILT_RANGE_EXT_RSTVAL : std_logic := '0';
  constant FILT_RANGE_BASIC_RSTVAL : std_logic := '0';
  constant FILT_C_FD_EXT_RSTVAL : std_logic := '0';

  ------------------------------------------------------------------------------
  -- FILTER_RAN_HIGH register
  --
  -- Higher threshold of the Range filter. Note that 29-bit value of range thres
  -- hold is not the same format as transmitted
  ------------------------------------------------------------------------------
  constant BIT_RAN_HIGH_VAL_L     : natural := 0;
  constant BIT_RAN_HIGH_VAL_H    : natural := 28;

  --FILTER_RAN_HIGH reset values
  constant BIT_RAN_HIGH_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_RAN_LOW register
  --
  -- Lower threshold of the Range filter. Note that 29-bit value of range thresh
  -- old is not the same format as transmitted and received identifier! In TX_DA
  -- TA_4 (transmitted identifier) BASE Identifier is at 11 LSB bits and Extensi
  -- on at bits 28-12. However, actual decimal value of the Identifier is that B
  -- ASE identifier is at MSB bits and 18 LSB bits is identifier extension. The 
  -- unsigned binary value of the identifier must be written into this register!
  --  Note that filter support is available by default but it can be left out fr
  -- om synthesis (to save logic) by setting "sup_ran=false". If the particular 
  -- filter is not supported, writes to this register have no effect and read wi
  -- ll return all zeroes.
  ------------------------------------------------------------------------------
  constant BIT_RAN_LOW_VAL_L      : natural := 0;
  constant BIT_RAN_LOW_VAL_H     : natural := 28;

  --FILTER_RAN_LOW reset values
  constant BIT_RAN_LOW_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_C_VAL register
  --
  -- Bit value for acceptance filters. Filters A, B, C are available. The identi
  -- fier format is the same as transmitted and
  ------------------------------------------------------------------------------
  constant BIT_VAL_C_VAL_L        : natural := 0;
  constant BIT_VAL_C_VAL_H       : natural := 28;

  --FILTER_C_VAL reset values
  constant BIT_VAL_C_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_C_MASK register
  --
  -- Bit mask for acceptance filters. Filters A, B, C are available. The identif
  -- ier format is the same as transmitted and
  ------------------------------------------------------------------------------
  constant BIT_MASK_C_VAL_L       : natural := 0;
  constant BIT_MASK_C_VAL_H      : natural := 28;

  --FILTER_C_MASK reset values
  constant BIT_MASK_C_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_B_VAL register
  --
  -- Bit value for acceptance filters. Filters A, B, C are available. The identi
  -- fier format is the same as transmitted and
  ------------------------------------------------------------------------------
  constant BIT_VAL_B_VAL_L        : natural := 0;
  constant BIT_VAL_B_VAL_H       : natural := 28;

  --FILTER_B_VAL reset values
  constant BIT_VAL_B_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_B_MASK register
  --
  -- Bit mask for acceptance filters. Filters A, B, C are available. The identif
  -- ier format is the same as transmitted and
  ------------------------------------------------------------------------------
  constant BIT_MASK_B_VAL_L       : natural := 0;
  constant BIT_MASK_B_VAL_H      : natural := 28;

  --FILTER_B_MASK reset values
  constant BIT_MASK_B_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- FILTER_A_MASK register
  --
  -- Bit mask for acceptance filters. Filters A, B, C are available. The identif
  -- ier format is the same as transmitted and received identifier format. BASE 
  -- Identifier is 11 LSB and Identifier extension are bits 28-12! Note that fil
  -- ter support is available by default but it can be left out from synthesis (
  -- to save logic) by setting "sup_fillt=false". If the particular filter is no
  -- t supported, writes to this register have no effect and read will return al
  -- l zeroes.
  ------------------------------------------------------------------------------
  constant BIT_MASK_A_VAL_L       : natural := 0;
  constant BIT_MASK_A_VAL_H      : natural := 28;

  --FILTER_A_MASK reset values
  constant BIT_MASK_A_VAL_RSTVAL : std_logic_vector(28 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- CTR_PRES register
  --
  -- Register for manipulation with error counters.
  ------------------------------------------------------------------------------
  constant CTR_PRES_VAL_L         : natural := 0;
  constant CTR_PRES_VAL_H         : natural := 8;
  constant PTX_IND                : natural := 9;
  constant PRX_IND               : natural := 10;
  constant ENORM_IND             : natural := 11;
  constant EFD_IND               : natural := 12;

  --CTR_PRES reset values
  constant CTR_PRES_VAL_RSTVAL : std_logic_vector(8 downto 0) := (OTHERS => '0');
  constant PTX_RSTVAL         : std_logic := '0';
  constant PRX_RSTVAL         : std_logic := '0';
  constant ENORM_RSTVAL       : std_logic := '0';
  constant EFD_RSTVAL         : std_logic := '0';

  ------------------------------------------------------------------------------
  -- ERR_FD register
  --
  ------------------------------------------------------------------------------
  constant ERR_FD_VAL_L          : natural := 16;
  constant ERR_FD_VAL_H          : natural := 31;

  --ERR_FD reset values
  constant ERR_FD_VAL_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- ERR_NORM register
  --
  -- Error counter for nominal Bit time
  ------------------------------------------------------------------------------
  constant ERR_NORM_VAL_L         : natural := 0;
  constant ERR_NORM_VAL_H        : natural := 15;

  --ERR_NORM reset values
  constant ERR_NORM_VAL_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- TXC register
  --
  -- Counter for transcieved frames to enable bus traffic measurement.
  ------------------------------------------------------------------------------
  constant TXC_VAL_L             : natural := 16;
  constant TXC_VAL_H             : natural := 31;

  --TXC reset values
  constant TXC_VAL_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');

  ------------------------------------------------------------------------------
  -- RXC register
  --
  -- Counter for received frames to enable bus traffic measurement.
  ------------------------------------------------------------------------------
  constant RXC_VAL_L              : natural := 0;
  constant RXC_VAL_H             : natural := 15;

  --RXC reset values
  constant RXC_VAL_RSTVAL : std_logic_vector(15 downto 0) := (OTHERS => '0');

  ----------------------------------------------------------------------------
  -- Address block: Control_Registers
  ----------------------------------------------------------------------------
  constant CONTROL_REGISTERS_BLOCK      : std_logic_vector(3 downto 0) := x"0";

  constant DEVICE_ID_ADR             : std_logic_vector(11 downto 0) := x"000";
  constant MODE_REG_ADR              : std_logic_vector(11 downto 0) := x"001";
  constant INTERRUPT_REG_ADR         : std_logic_vector(11 downto 0) := x"002";
  constant TIMING_REG_ADR            : std_logic_vector(11 downto 0) := x"003";
  constant ARB_ERROR_PRESC_ADR       : std_logic_vector(11 downto 0) := x"004";
  constant ERROR_TH_ADR              : std_logic_vector(11 downto 0) := x"005";
  constant ERROR_COUNTERS_ADR        : std_logic_vector(11 downto 0) := x"006";
  constant ERROR_COUNTERS_SPEC_ADR   : std_logic_vector(11 downto 0) := x"007";
  constant CTR_PRES_ADR              : std_logic_vector(11 downto 0) := x"008";
  constant FILTER_A_VAL_ADR          : std_logic_vector(11 downto 0) := x"009";
  constant FILTER_A_MASK_ADR         : std_logic_vector(11 downto 0) := x"00A";
  constant FILTER_B_VAL_ADR          : std_logic_vector(11 downto 0) := x"00B";
  constant FILTER_B_MASK_ADR         : std_logic_vector(11 downto 0) := x"00C";
  constant FILTER_C_VAL_ADR          : std_logic_vector(11 downto 0) := x"00D";
  constant FILTER_C_MASK_ADR         : std_logic_vector(11 downto 0) := x"00E";
  constant FILTER_RAN_LOW_ADR        : std_logic_vector(11 downto 0) := x"00F";
  constant FILTER_RAN_HIGH_ADR       : std_logic_vector(11 downto 0) := x"010";
  constant FILTER_CONTROL_ADR        : std_logic_vector(11 downto 0) := x"011";
  constant RX_INFO_1_ADR             : std_logic_vector(11 downto 0) := x"012";
  constant RX_INFO_2_ADR             : std_logic_vector(11 downto 0) := x"013";
  constant RX_DATA_ADR               : std_logic_vector(11 downto 0) := x"014";
  constant TRV_DELAY_ADR             : std_logic_vector(11 downto 0) := x"015";
  constant TX_STATUS_ADR             : std_logic_vector(11 downto 0) := x"016";
  constant TX_SETTINGS_ADR           : std_logic_vector(11 downto 0) := x"017";
  constant ERR_CAPT_ADR              : std_logic_vector(11 downto 0) := x"018";
  constant RX_COUNTER_ADR            : std_logic_vector(11 downto 0) := x"02B";
  constant TX_COUNTER_ADR            : std_logic_vector(11 downto 0) := x"02C";
  constant LOG_TRIG_CONFIG_ADR       : std_logic_vector(11 downto 0) := x"02E";
  constant LOG_CAPT_CONFIG_ADR       : std_logic_vector(11 downto 0) := x"030";
  constant LOG_STATUS_ADR            : std_logic_vector(11 downto 0) := x"031";
  constant LOG_CMD_ADR               : std_logic_vector(11 downto 0) := x"032";
  constant LOG_CAPT_EVENT_1_ADR      : std_logic_vector(11 downto 0) := x"033";
  constant LOG_CAPT_EVENT_2_ADR      : std_logic_vector(11 downto 0) := x"034";
  constant DEBUG_REG_ADR             : std_logic_vector(11 downto 0) := x"035";
  constant YOLO_REG_ADR              : std_logic_vector(11 downto 0) := x"036";


  ----------------------------------------------------------------------------
  -- Address block: TX_Buffer
  ----------------------------------------------------------------------------
  constant TX_BUFFER_BLOCK              : std_logic_vector(3 downto 0) := x"1";

  constant TX_DATA_1_ADR             : std_logic_vector(11 downto 0) := x"100";
  constant TX_DATA_2_ADR             : std_logic_vector(11 downto 0) := x"101";
  constant TX_DATA_3_ADR             : std_logic_vector(11 downto 0) := x"102";
  constant TX_DATA_4_ADR             : std_logic_vector(11 downto 0) := x"103";
  constant TX_DATA_5_ADR             : std_logic_vector(11 downto 0) := x"104";
  constant TX_DATA_6_ADR             : std_logic_vector(11 downto 0) := x"105";
  constant TX_DATA_7_ADR             : std_logic_vector(11 downto 0) := x"106";
  constant TX_DATA_8_ADR             : std_logic_vector(11 downto 0) := x"107";
  constant TX_DATA_9_ADR             : std_logic_vector(11 downto 0) := x"108";
  constant TX_DATA_10_ADR            : std_logic_vector(11 downto 0) := x"109";
  constant TX_DATA_11_ADR            : std_logic_vector(11 downto 0) := x"10A";
  constant TX_DATA_12_ADR            : std_logic_vector(11 downto 0) := x"10B";
  constant TX_DATA_13_ADR            : std_logic_vector(11 downto 0) := x"10C";
  constant TX_DATA_14_ADR            : std_logic_vector(11 downto 0) := x"10D";
  constant TX_DATA_15_ADR            : std_logic_vector(11 downto 0) := x"10E";
  constant TX_DATA_16_ADR            : std_logic_vector(11 downto 0) := x"10F";
  constant TX_DATA_17_ADR            : std_logic_vector(11 downto 0) := x"110";
  constant TX_DATA_18_ADR            : std_logic_vector(11 downto 0) := x"111";
  constant TX_DATA_19_ADR            : std_logic_vector(11 downto 0) := x"112";
  constant TX_DATA_20_ADR            : std_logic_vector(11 downto 0) := x"113";


end package;