--------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core
-- Copyright (C) 2015-2018
-- 
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <jerabma7@fel.cvut.cz>
-- 
-- Project advisors: 
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
-- 
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy 
-- of this VHDL component and associated documentation files (the "Component"), 
-- to deal in the Component without restriction, including without limitation 
-- the rights to use, copy, modify, merge, publish, distribute, sublicense, 
-- and/or sell copies of the Component, and to permit persons to whom the 
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in 
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR 
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY, 
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE 
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER 
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS 
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents. 
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN 
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------


configuration tbconf_{{test}} of vunittb_wrapper is
for tb
    for i_test : CAN_test use entity work.CAN_test({{test}}); end for;
end for;
end configuration;
-- -----------------------------------------------------------------------------
{% endfor %}

-- Entities
{% for test in tests %}

library work;
use work.CANtestLib.all;
library vunit_lib;
context vunit_lib.vunit_context;

entity tb_{{test}} is generic (
    runner_cfg : string := runner_cfg_default;
    iterations : natural := 1;
    log_level  : log_lvl_type := info_l;
    error_beh  : err_beh_type := quit;
    error_tol  : natural := 0;
    timeout    : string := "0 ms";
    seed       : natural := 0
); end entity;
architecture tb of tb_{{test}} is
    component vunittb_wrapper is generic (
        nested_runner_cfg : string;
        iterations : natural;
        log_level  : log_lvl_type;
        error_beh  : err_beh_type;
        error_tol  : natural;
        timeout    : string;
        seed       : natural
    ); end component;
    for all:vunittb_wrapper use configuration work.tbconf_{{test}};
begin
    tb:vunittb_wrapper generic map(
        nested_runner_cfg => runner_cfg,
        iterations        => iterations,
        log_level         => log_level,
        error_beh         => error_beh,
        error_tol         => error_tol,
        timeout           => timeout,
        seed              => seed);
end architecture;
-- -----------------------------------------------------------------------------
{% endfor %}
