--------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core 
-- Copyright (C) 2021-present Ondrej Ille
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to use, copy, modify, merge, publish, distribute the Component for
-- educational, research, evaluation, self-interest purposes. Using the
-- Component for commercial purposes is forbidden unless previously agreed with
-- Copyright holder.
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
-- -------------------------------------------------------------------------------
-- 
-- CTU CAN FD IP Core 
-- Copyright (C) 2015-2020 MIT License
-- 
-- Authors:
--     Ondrej Ille <ondrej.ille@gmail.com>
--     Martin Jerabek <martin.jerabek01@gmail.com>
-- 
-- Project advisors: 
-- 	Jiri Novak <jnovak@fel.cvut.cz>
-- 	Pavel Pisa <pisa@cmp.felk.cvut.cz>
-- 
-- Department of Measurement         (http://meas.fel.cvut.cz/)
-- Faculty of Electrical Engineering (http://www.fel.cvut.cz)
-- Czech Technical University        (http://www.cvut.cz/)
-- 
-- Permission is hereby granted, free of charge, to any person obtaining a copy
-- of this VHDL component and associated documentation files (the "Component"),
-- to deal in the Component without restriction, including without limitation
-- the rights to use, copy, modify, merge, publish, distribute, sublicense,
-- and/or sell copies of the Component, and to permit persons to whom the
-- Component is furnished to do so, subject to the following conditions:
-- 
-- The above copyright notice and this permission notice shall be included in
-- all copies or substantial portions of the Component.
-- 
-- THE COMPONENT IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
-- IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
-- FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
-- AUTHORS OR COPYRIGHTHOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
-- LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
-- FROM, OUT OF OR IN CONNECTION WITH THE COMPONENT OR THE USE OR OTHER DEALINGS
-- IN THE COMPONENT.
-- 
-- The CAN protocol is developed by Robert Bosch GmbH and protected by patents.
-- Anybody who wants to implement this IP core on silicon has to obtain a CAN
-- protocol license from Bosch.
-- 
--------------------------------------------------------------------------------

--------------------------------------------------------------------------------
-- @TestInfoStart
--
-- @Purpose:
--  STATUS[TXNF] feature test.
--
-- @Verifies:
--  @1. When no TXT Buffer is in Empty state, STATUS[TXNF] is not set.
--  @2. When at least on TXT Buffer is in Empty state STATUS[TXNF] is set.
--
-- @Test sequence:
--  @1. Set BMM mode in Node 1. Check that STATUS[TXNF] is set (all TXT Buffers
--      should be empty).
--  @2. Issue Set ready consecutively to all TXT Buffers. Check that STATUS[TXNF]
--      is set before last buffer. Check that after last buffer STATUS[TXNF] is
--      not set.
--  @3. Check that all TXT Buffers are Failed now. Move always single buffer to
--      empty and check that STATUS[TXNF] is set. Move this buffer to Failed again
--      and check that STATUS[TXNF] is not set. Repeat with each TXT Buffer.
--
-- @TestInfoEnd
--------------------------------------------------------------------------------
-- Revision History:
--    31.10.2019   Created file
--------------------------------------------------------------------------------

Library ctu_can_fd_tb;
context ctu_can_fd_tb.ctu_can_synth_context;
context ctu_can_fd_tb.ctu_can_test_context;

use ctu_can_fd_tb.pkg_feature_exec_dispath.all;

package status_txnf_feature is
    procedure status_txnf_feature_exec(
        signal      so              : out    feature_signal_outputs_t;
        signal      rand_ctr        : inout  natural range 0 to RAND_POOL_SIZE;
        signal      iout            : in     instance_outputs_arr_t;
        signal      mem_bus         : inout  mem_bus_arr_t;
        signal      bus_level       : in     std_logic
    );
end package;


package body status_txnf_feature is
    procedure status_txnf_feature_exec(
        signal      so              : out    feature_signal_outputs_t;
        signal      rand_ctr        : inout  natural range 0 to RAND_POOL_SIZE;
        signal      iout            : in     instance_outputs_arr_t;
        signal      mem_bus         : inout  mem_bus_arr_t;
        signal      bus_level       : in     std_logic
    ) is
        variable ID_1               :     natural := 1;
        variable ID_2               :     natural := 2;

        -- Generated frames
        variable frame_1            :     SW_CAN_frame_type;

        -- Node status
        variable stat_1             :     SW_status;
        
        variable txt_buf_state      :     SW_TXT_Buffer_state_type;
        variable mode_1             :     SW_mode;
    begin

        -----------------------------------------------------------------------
        -- @1. Set BMM mode in Node 1. Check that STATUS[TXNF] is set (all TXT
        --    Buffers should be empty).
        -----------------------------------------------------------------------
        info("Step 1");
        mode_1.bus_monitoring := true;
        set_core_mode(mode_1, ID_1, mem_bus(1));

        get_controller_status(stat_1, ID_1, mem_bus(1));
        check(stat_1.tx_buffer_empty, "STATUS[TXNF] set!");

        -----------------------------------------------------------------------
        -- @2. Issue Set ready consecutively to all TXT Buffers. Check that
        --     STATUS[TXNF] is set before last buffer. Check that after last
        --     buffer STATUS[TXNF] is not set.
        -----------------------------------------------------------------------
        for i in 1 to C_TXT_BUFFER_COUNT loop
            send_TXT_buf_cmd(buf_set_ready, i, ID_1, mem_bus(1));

            get_controller_status(stat_1, ID_1, mem_bus(1));

            if (i = C_TXT_BUFFER_COUNT) then
                check_false(stat_1.tx_buffer_empty,
                    "STATUS[TXNF] not set after last TXT Buffer");
            else
                check(stat_1.tx_buffer_empty,
                    "STATUS[TXNF] set before last TXT Buffer");
            end if;
        end loop;

        -----------------------------------------------------------------------
        -- @3. Check that all TXT Buffers are Failed now. Move always single
        --    buffer to empty and check that STATUS[TXNF] is set. Move this
        --    buffer to Failed again and check that STATUS[TXNF] is not set.
        --    Repeat with each TXT Buffer.
        -----------------------------------------------------------------------
        info("Step 3");
        for i in 1 to C_TXT_BUFFER_COUNT loop
            get_tx_buf_state(i, txt_buf_state, ID_1, mem_bus(1));
            check(txt_buf_state = buf_failed, "TXT Buffer: " &
                integer'image(i) & " failed!");
        end loop;

        for i in 1 to C_TXT_BUFFER_COUNT loop
            send_TXT_buf_cmd(buf_set_empty, i, ID_1, mem_bus(1));
            
            get_controller_status(stat_1, ID_1, mem_bus(1));
            check(stat_1.tx_buffer_empty, "STATUS[TXNF] set!");
            
            send_TXT_buf_cmd(buf_set_ready, i, ID_1, mem_bus(1));
            
            get_controller_status(stat_1, ID_1, mem_bus(1));
            check_false(stat_1.tx_buffer_empty, "STATUS[TXNF] not set!");
            
            get_tx_buf_state(i, txt_buf_state, ID_1, mem_bus(1));
            check(txt_buf_state = buf_failed, "TXT Buffer: " &
                integer'image(i) & " ready!");
        end loop;
        
        wait for 100 ns;

  end procedure;

end package body;
